--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.9 Beta-4 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Sun Dec 31 19:10:45 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_basic_kernal is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_basic_kernal;

architecture Behavioral of Gowin_pROM_basic_kernal is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"39556CEAE29F59569B269A2452FA5E4BE8F66139EE05AF5456BC890C64A7CF5E",
            INIT_RAM_01 => X"D132A248E13A3129494AAD2D998C21E85714F9C1E8E9692B548A459F57B2C649",
            INIT_RAM_02 => X"4ECB54AA652BEA68E691EB2745B23A94DE4F169CE689BCCC5268CC4B3A39E52F",
            INIT_RAM_03 => X"9052C5215529839D1804AF77F46F80E2564448FEA910110154EABA6A9A8A74CB",
            INIT_RAM_04 => X"EE0E42A2A949E2EBEDEBFC2B6D820A248C990960364CB67DA20B800D4190C001",
            INIT_RAM_05 => X"8D03A62DB311F9631102291B3A1641C608154370589D09226498C87519EB3250",
            INIT_RAM_06 => X"FC773A00F32175B9A191896B07AF8A800919999E90AEBD98B30664796719EE10",
            INIT_RAM_07 => X"265C93290A5694490C121B21446A4A9B5D992C9C9361A996C1410A6ABA49B31C",
            INIT_RAM_08 => X"A4C96450B479ABE231496BB681364BDA0A44339D41455866609161A3C12AE0E4",
            INIT_RAM_09 => X"05414448211ED3204232935943B1EA809BFD00396159A612B5AED4A422721010",
            INIT_RAM_0A => X"503C4879AD9D16D96287313A58244D306B5A293072904DB046A949883B842122",
            INIT_RAM_0B => X"C6A58461D7BB32D4A272498A4B4A4988E24E4A2E19916E6CDC56C8008C102C2F",
            INIT_RAM_0C => X"341BB151A2249685044A52673A6514A44994ECE68AA51B5C518428239345A4A6",
            INIT_RAM_0D => X"81A227577165DFBBB2D5B008112A1229469F6B7F71511BD22908A1A812B1555A",
            INIT_RAM_0E => X"25C1A65ED7E89893332636506E594B63D596592D320CB2D1840CDA3183710142",
            INIT_RAM_0F => X"47FDD0B07F4502059940484918081C44254530890408842022994A7A8EA84A52",
            INIT_RAM_10 => X"79861869422F51B3C4D25A444B2C4040862229444278CC81318B511AED37EB7F",
            INIT_RAM_11 => X"FABA85A320CA8573CE89380947B1A17B6D9D786992B4999C1CAA935C8DD8BCB2",
            INIT_RAM_12 => X"3C877C3A73D452A13024EC86999301B1C1A5F0082CE4C8139B1A6CA166759429",
            INIT_RAM_13 => X"45ED2156816C92B2513290260130AF416A98910006F9C676B202B92B050692B0",
            INIT_RAM_14 => X"8DA02840FAEA80124888F49933526438110198C44444652594674A5C03326996",
            INIT_RAM_15 => X"0AFE6588120514853612A17084F4A88922E27E6D6127F69933321986C3019D90",
            INIT_RAM_16 => X"021661E98201E5441110A6703C1A0833320060484A962D9171715693D5DC79C5",
            INIT_RAM_17 => X"7CC5A20909224A94050A8A091084210A401E418577881688D7CD6010A025010E",
            INIT_RAM_18 => X"4E8A41410069DE977A57455495810384187048187AE856350D22C46991316C95",
            INIT_RAM_19 => X"3AF109405A9087661008A88483050412810103BFBBFBAE88823FB044715FD5FD",
            INIT_RAM_1A => X"00A5020222D3AB4235BD2BAAD2B490110AFEAFE8B582B4AD3BAA50B852AC4EB5",
            INIT_RAM_1B => X"50E5D394E422080D2AB4AD257AFAA3100715FD5FC0110C3450050184BCA04906",
            INIT_RAM_1C => X"E901BA3F4888711450C733A11AC4D74A352B4282480B3AD354CCDC34588A2116",
            INIT_RAM_1D => X"8194A5E0D321332C9CCC520890CA2D402441122E05021CD5920223133918CAC8",
            INIT_RAM_1E => X"B5D925FE481A44E003A9927941B80035FED7EC264334252CE5C910200AC14F8B",
            INIT_RAM_1F => X"0A5161138C2DE03C9D30C06124844C0564B0000000001C1D8FC1D0C941009AB2",
            INIT_RAM_20 => X"81096BA9B1B21070D6B45291891042146B18302FC60D0E19354C4B2EE6B604E9",
            INIT_RAM_21 => X"90248110D1956D2896124A0EABC932CE26C4C56A651D3504D5CBC04102D84844",
            INIT_RAM_22 => X"ED9884E74C21586012C472218ECA8815A060C21D0A0130022B003428B32480A0",
            INIT_RAM_23 => X"A69D7C74393B9C6A98948980432124036063840D61E3071F5201B29D36E44EEF",
            INIT_RAM_24 => X"56F7F58965790B801D9190191300F057C01B8D3CA5715388395B860C1608B0A0",
            INIT_RAM_25 => X"E8488F2849A2B0083224E6D7906C3089C1A2C2063E0944975A52D3B76C448900",
            INIT_RAM_26 => X"D0497ADBA8051A277C80010800925D131C3E5056B024012BFA421D28590049C8",
            INIT_RAM_27 => X"A87A615A94F0803103096201492E5E2A2CED36D845B015086622AE5CA1950440",
            INIT_RAM_28 => X"789966AD2800302015E005680441031424910C61143D1A18B20D300CED36D858",
            INIT_RAM_29 => X"13F96FA84DDA6781052D95A8AC144CB202002B05960DF78687988AC236CAE456",
            INIT_RAM_2A => X"7703234E408944366780D82BFA918680D7E2380E143C35AADA985DF6E0D03409",
            INIT_RAM_2B => X"0EF4A5CD1C479F5B877812E68E23CFAC361BF2285330DB1C31020A8081421266",
            INIT_RAM_2C => X"0000FF5528040C0001FCB6B9724710EEFD0DE73641CCC99E5DF113A8F746D477",
            INIT_RAM_2D => X"DD681A21049485AF56032085B7B4ABD04A150B744A522428482B64C689009200",
            INIT_RAM_2E => X"119F70C5DB280A7021005AAD5EAB57A1100A1690B7482846C14B69EF92D24826",
            INIT_RAM_2F => X"02C46D9681CB10CDE2140E8F5D4B160800270B3408030404F3102140F3106163",
            INIT_RAM_30 => X"C64D2271B9255F25F6F4261210969FB63733886A86207099C0538CF9B3A91A00",
            INIT_RAM_31 => X"C33723B0661068FFCF4629300600384CC8C076C6BD812A04C899D78DB555EB72",
            INIT_RAM_32 => X"D8002580296422371B04A546260981A9700C81AF4ED6C0C21E16391963B5B02A",
            INIT_RAM_33 => X"B0F139E2A4610B1528C14483733536EB4635EED1402D21A6A912B6B587028DB6",
            INIT_RAM_34 => X"ACBAD71A055BCEDD2AAF4AF0858A65302602E4027CC825FA45088039A5F91C09",
            INIT_RAM_35 => X"BEBD31F51A384985ABC1A06D8853C0800C0769185B4200112DA4868810442024",
            INIT_RAM_36 => X"58C5E1224C112141B20D7D0406D5989DC5509A00584CFC6A4845B22DE61B8AD2",
            INIT_RAM_37 => X"D97D76947664A94A5A299560B41644AA29C3400648DAC2E51C8B811311196596",
            INIT_RAM_38 => X"D866852000860B328A8C4456400C0862BA20920814AF690150227001A0326078",
            INIT_RAM_39 => X"4B16076CAC8E3172924441D4D541529572C63BE4A4022CD123DEF0F932CF2802",
            INIT_RAM_3A => X"94B7BAD0EEB4F1E6014D81068BA1B209D2B639BFE088C1E548B86400D802F9C0",
            INIT_RAM_3B => X"0673A8C116F20E010F3395A6601F4003C0644AFE529B23A9CE27068E4144080A",
            INIT_RAM_3C => X"3698080903D4DD057DE0C0CF0D602C22BC6609DB24FA0C19A3635B0014522128",
            INIT_RAM_3D => X"171A7C9C2FF7B80C8EE94F7AA14A80083DFE89440249D39BC1914BDB890549F8",
            INIT_RAM_3E => X"150703244C6AE6380EC026A2009A1401A2784D80050DF04020804106571A72A1",
            INIT_RAM_3F => X"8624CA4886124924C169364905B09A6D074BF1DC64534012CC3C15418C822AF2"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"9A2AA43A9C6ED6B6040A201E87D67BD0EAE23BA5BA02D0ADF704544440E48ABE",
            INIT_RAM_01 => X"0813108D519459864C321891980A45C5644978CEE7B2E75D170BC94B669A8EAA",
            INIT_RAM_02 => X"06C0E01E66A88050434B50C423D1409930C76C204018DC4588BC4434941010B6",
            INIT_RAM_03 => X"2AB902108752892A401991290A80049CA188F06EFAABEBFFEA444125734C89CD",
            INIT_RAM_04 => X"502295C13A28495009045068282F2AC686A52D183489A25ADE222041AB0A8056",
            INIT_RAM_05 => X"41E1228428249040243A000022A2055239960809170A31408510504144241014",
            INIT_RAM_06 => X"AAB4002026615014049503222515040E344141160D012900A64404414C32B141",
            INIT_RAM_07 => X"00D01A29D4A114AA20D40051250306AAAA4301090B074C00D21218CAAB60E610",
            INIT_RAM_08 => X"429204498EA1045661711002C00092D2924082A15761405103A044008308A504",
            INIT_RAM_09 => X"883A1016290001280905A841310A107E0454A909608034108068022804D81ADD",
            INIT_RAM_0A => X"1088885A2C11C2D1085512281206C1A60000600C40020401142825485895A848",
            INIT_RAM_0B => X"9495504AC511A6A5365978CB442578C8B2A3024A411008405490D11CAD954303",
            INIT_RAM_0C => X"160AA14902842508D21014455220A41600A05544600572501C000B32A8460246",
            INIT_RAM_0D => X"90205A9150A4004A800D847ED628082019D0940504114438106B3428049D30F1",
            INIT_RAM_0E => X"002DA24484288C8154454D5A2A494830A80482A112412011383406020117DED6",
            INIT_RAM_0F => X"42285080B18993204A2C4AE01A2904E4A0412420450214002044821100040B54",
            INIT_RAM_10 => X"4504E0081A908080A252C85AC90108030559BA05D2A4011C1664050554254221",
            INIT_RAM_11 => X"040148104010A4001048080004610252490A4040802541101488885101002824",
            INIT_RAM_12 => X"A0482910AA09B00C812200E9950400E13D490C01A8846B713255080233283500",
            INIT_RAM_13 => X"89414830824835820DA2C8E2034B022D0982568B8810A40460F506B4932104AA",
            INIT_RAM_14 => X"0936300944092E185061202822544F8B0231080888884921224294942204D520",
            INIT_RAM_15 => X"D48BB8C88AA265085280FA890C081131DA29292041D9522E46CA0CC42A4C1404",
            INIT_RAM_16 => X"4400C15102CD45442621A81380044B26202C53060B0408B00A0E064682A10287",
            INIT_RAM_17 => X"016992E4080023C9F36AC11094C830BB6400100C014274D20168451D41802404",
            INIT_RAM_18 => X"90002AEFD82A0522400A10504400C151020ECA01155450083905C0EC00300005",
            INIT_RAM_19 => X"40894980421BA73E005F56404011440ADDCCC90411555515F98285EA8AAA8000",
            INIT_RAM_1A => X"0095B42120A5280004024554A108A52BF554000055B528420146D40440800624",
            INIT_RAM_1B => X"A10AA52105A90C82452842290055270FE32AA800157AC08100151433802A6DB0",
            INIT_RAM_1C => X"2A6014A02508002B2010C14840A80240A0401410035081A6242B0094C121A241",
            INIT_RAM_1D => X"209209141903CCA0EF58843340149A80120CD208F478A15621026228A905488C",
            INIT_RAM_1E => X"0AAA380181708088096129544151A85AB44081042A455A5A88280E9D48A90140",
            INIT_RAM_1F => X"0A0940266517FB162A8A9091A48854310681FFFFFFF80D1D9FE1D0D051C00020",
            INIT_RAM_20 => X"BB0D00431E4A2818912825178921030500448E08D1084B42204444401084240A",
            INIT_RAM_21 => X"CB1648B60301622932CB555492CD15466A8708025219AC06B190D84580986C90",
            INIT_RAM_22 => X"85B607BC8C528C48F465522A951010A5006E0289796D8D9B083984DD21210436",
            INIT_RAM_23 => X"494828D92288D220380454ECEB212C5A203F19CAC07706ABD20882AC1024BA95",
            INIT_RAM_24 => X"004004025914C051772300DA10F6A934DE0868AAAC5F63CC0032C408DC0CE0E3",
            INIT_RAM_25 => X"2B964968F12C583268E5C30A400908210300BA2A4A80104025A989628058B821",
            INIT_RAM_26 => X"8183002017D46AD5468218DBB2588022A8A35748113210AE8A128A81C1604800",
            INIT_RAM_27 => X"A80224448AA8B020E0C01A060921555A4B04240241A48D3A5400225403103876",
            INIT_RAM_28 => X"27D20333A1C45B8D455B514786EA3050D48C2B4D008820502EE3039B05240200",
            INIT_RAM_29 => X"290044440A08121A988AA68008A0A901BD44586024F000805428100029402000",
            INIT_RAM_2A => X"445AB112C04B05484028011500888810311000410BEA587E010C0A8524250141",
            INIT_RAM_2B => X"AB21C79254E8CD83559C63C92A7466C03D2C4D1C204B140B6A78D0858BD48000",
            INIT_RAM_2C => X"0000596636040C0001B6F8B9ED9D3ABAFFD25042300510AF1651BC94DB115946",
            INIT_RAM_2D => X"900600040522C004011201280420410F9A8340035294A840DB001420D1A00000",
            INIT_RAM_2E => X"420A90545B202A20925A000008000200D10480240026122802501908A40693D0",
            INIT_RAM_2F => X"4210EC66241842011A4321A8012006CA8C0001840D084C5D0843B46708424008",
            INIT_RAM_30 => X"052000436076657994A0324A134D811155018504841CD702D9FAC56AD41E6104",
            INIT_RAM_31 => X"C8500580E0185102B2C0114006040C2006C600B15400002808D00316CA9AB124",
            INIT_RAM_32 => X"200D8479002141621180E1444E29A22402A8820A5696D15040E4BC8155A5A490",
            INIT_RAM_33 => X"20B0000415048904226100AD108C10EA156A010753ADA41A855809620858126D",
            INIT_RAM_34 => X"A8068A3632C814048A0B5050E8A3212AA20042AA240512A2E059C3CC9A2B8328",
            INIT_RAM_35 => X"822D5A0368A14D04A2442C1CA40A85DE98004C12D62862250104328EE408299D",
            INIT_RAM_36 => X"814500C1820012D00D68823368441801080235C8822040810835010C03001692",
            INIT_RAM_37 => X"4A229404D40129100028A942AC4802388011C0410D0A02208185218141004804",
            INIT_RAM_38 => X"0281401200A4160A2CC86A845E8BC01404440E842044208002081420A903010A",
            INIT_RAM_39 => X"C4E0A28020052F11490203032C020E0428010458414012025010A10A02AA1044",
            INIT_RAM_3A => X"AE0A508B94214A0C363410104A911540DA04215051829C05910C2A813B858D2F",
            INIT_RAM_3B => X"2A050451B2858360255105303700A49A8802218960A011040541110D501184E2",
            INIT_RAM_3C => X"30098B2CCA200002C450480240040517A01400888419451E624A50613626EB1B",
            INIT_RAM_3D => X"1D840402C44A1396D4920014843114700811205C89100F65EEFE09428C231924",
            INIT_RAM_3E => X"BD26268060C9035081008B282908D5DB1409040D148021435D64F3C80030C50C",
            INIT_RAM_3F => X"9DC21A69205A69A6130090D34884402DC81006048410224000C0B4F8C5C31E02"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"2BA7973B6B976ADFEAE9A5B7DCBE5000FBBF547194BA1479505510145C578041",
            INIT_RAM_01 => X"EB77D69FA3A7FBB75DBAD695DEE9F816BB6B11F82A46DDDA6FA1E3FDB4653D86",
            INIT_RAM_02 => X"6CE76ADF764529A57A83140ED024FD3F9EDFDD69795BADD5718DD56BA75ED6B0",
            INIT_RAM_03 => X"A02800915229029D2C008B14A44080226A4848B151501101144015B4F5DFFB9C",
            INIT_RAM_04 => X"AE0C83441161E3DFE9EBB1460B260161822814121404932D6081AC0561806349",
            INIT_RAM_05 => X"08A0062D308400A121091A88AB862547967C03404A04080A02ED9048FAB7E10E",
            INIT_RAM_06 => X"EE14998EE22459F5E4044200A36C8E00312BFEBE8D9E1008A214C0594E699519",
            INIT_RAM_07 => X"44405F028A4208003E0A8132410015585B9B4484880120924242094B29B9E210",
            INIT_RAM_08 => X"A24925E620688A76D9286E80E022490394405D5F993A01ABF158428C47402C32",
            INIT_RAM_09 => X"64A13A56A44631404337850467FFEFA5C3F5E1407585372004EA060120FA9908",
            INIT_RAM_0A => X"308A0848950910036BD142020082D59A00004508EBA0FDF1F32B8F10177828A2",
            INIT_RAM_0B => X"5250C4A8D21C863013293AC1C1013AC0117D5726ABD4295A0944440D80442502",
            INIT_RAM_0C => X"B3A9018ED800862102FA0BBAACA03944C05564762130A10D115205DD551A9168",
            INIT_RAM_0D => X"51A026E745D19E0080C801147D035B0200E94A5713012E40721C82809935D770",
            INIT_RAM_0E => X"5269C991B5A00B80B00144222A828309FDB2491C422496E0943DBC00016289D2",
            INIT_RAM_0F => X"25F749BAE709C30D9B68401FFA809BEE341589116F2E5E82B25FF866066A5C20",
            INIT_RAM_10 => X"59CEFA10580FC123AA00021E500F0201BC2028A5C2E604F9EAEF0A02D90BB95D",
            INIT_RAM_11 => X"73888D8360DF4840DEC1E8050F138472490B58E50A22ABBD45082F4408442CA6",
            INIT_RAM_12 => X"AD851872634CA0945804665551000C20A16172446A559E931A57681977EDB240",
            INIT_RAM_13 => X"8D8FE135C12CB1B04887304238B8E56C630882C006319656908639174C82BBA2",
            INIT_RAM_14 => X"35363CF8AABC8E3E04A17201BA4AEE15CBE118C888882541B4658C4A422471B6",
            INIT_RAM_15 => X"8A77D5CE91AC0001061951600050A000BC65514D72BED6B5075F35C66B07E8C2",
            INIT_RAM_16 => X"A0304199C958A0D8000117F33C10052222C8FA2CDEA42DA3762A5A5D45ECBBC2",
            INIT_RAM_17 => X"0DFDA15610446174AAAC873101202190C01A418D674004DA07784B88A1170084",
            INIT_RAM_18 => X"DA40EFBA8821428D1E9E00585424617A4A26B140BFDA701618018843B2336FF9",
            INIT_RAM_19 => X"48921100B581281C0235546440AABAF788D9CB3DF6CB3D9F519290BE8D557FFD",
            INIT_RAM_1A => X"82958019B2B7912A949427F84632542BFBEEEBA008D2118C2BE2222C40001204",
            INIT_RAM_1B => X"F221B08C72C58B1426118C95EEBBF990219557FFC52FC2107DE28A4294491181",
            INIT_RAM_1C => X"A181EA7D07B012153110130C0D8CE61C182427447B3AF89118098914890B4216",
            INIT_RAM_1D => X"00E21D460F40AB007BF5C01863065FF32E019B8CC4683D9F713068028815022E",
            INIT_RAM_1E => X"00002084C160809AA1352B50E1140A3973CF8C1422483C0A01905AB1120A470A",
            INIT_RAM_1F => X"30114007C2EB9F503B90C080B10B5A22208C000000061D0C0FC3C0D151000021",
            INIT_RAM_20 => X"E0C122E6EBBA00400E10C24B0A20CB24A228541C4A49082830560F156007903B",
            INIT_RAM_21 => X"A8044012018244083CD517C3EAC650C6A6DAA48A1E8CDB336CD0CC6596F84A0D",
            INIT_RAM_22 => X"84AB84846649C04882025820CC9898019B2CB20EB325140A0110841C3161803A",
            INIT_RAM_23 => X"1B151026D0F0240F18040146114FC111300372C4771BC9E49C0080245070C8F6",
            INIT_RAM_24 => X"5A97D4C40FB482805901008E3B02035F8013A600A1E7DC751B4B51358835E373",
            INIT_RAM_25 => X"A8FE020C7DA3F83B3234F644F192F82508817D021800201F88E26233243E7808",
            INIT_RAM_26 => X"459038C897C46C253A0011C1E21833022C3B030C9390B83EC440151D8E91401C",
            INIT_RAM_27 => X"A60EAC9508A63A18CBC11D16642B061CE18580012164AE3745004B9A818FB436",
            INIT_RAM_28 => X"679B6C3BF8C2330D04C34121D3E9F900DE0FA3CE802C8B0C1EE393D18480016A",
            INIT_RAM_29 => X"122D61FA42286431C4199C80FE980DB77314316DB6F451820C8A0F6027D54AAB",
            INIT_RAM_2A => X"444681696A880236152168B660AD4601D3320A028DB1783DEB38C15012C10221",
            INIT_RAM_2B => X"1B92734315B5283E0DC339A18ADA94EF407394064319C35B38EA6F66688E7145",
            INIT_RAM_2C => X"000085F84606080001BEF79DD0CD6DCBFFE4D012398901A87736F8A5B4A1CA74",
            INIT_RAM_2D => X"B52E1A2D613685AD56188503FE7AE950D8970B7310841D429B294906788D4800",
            INIT_RAM_2E => X"953DD0419B00F48021205AA55AA956A3C32E16F0B70F1A52CA47FB9C26CFC834",
            INIT_RAM_2F => X"00E3F974B29C56E1FE4E150FC972E6C0BF2749AC4C038D195B95F0F75B9420DB",
            INIT_RAM_30 => X"124E074AA5360A25B0A4000003A30B010501A52206206282D072613A618C0A00",
            INIT_RAM_31 => X"C1150180575D08ED9DA526E00410047CC6A5742BA88943AE40915DBFC9DA75F9",
            INIT_RAM_32 => X"43290D8619A30FDD9910E0502205C50D388801038AA2F2C74C14D10C12A8B818",
            INIT_RAM_33 => X"82F9307296255DD9459D46045BB145595015A25683C5448E1C22169483120D10",
            INIT_RAM_34 => X"48B5FD1C07998A4CA3828A27448D2724B230E34A5424A4C840044894A4491DED",
            INIT_RAM_35 => X"D20A2555E4116816AB55BD587EF147CC0C144C105B6240783837261CEE089029",
            INIT_RAM_36 => X"21E522A54452DB02D569112325419C9965098B6848684E475025354FED11CE54",
            INIT_RAM_37 => X"471C60ABA610701111088145061200A325169C23484820E38B8BA1011984DB69",
            INIT_RAM_38 => X"F470C032E12420C5DD335804000FE0FE9480B6C415AD4BDD02111820813A4B68",
            INIT_RAM_39 => X"0120A5270E621060A3065852B96158A3629F2BAF9D1CE707F1F9ED78E00A31DE",
            INIT_RAM_3A => X"0C977A59DE94CC8FF90845A02020802AFCB02098E8CE88A5C4042204A801C864",
            INIT_RAM_3B => X"C62295F326A3846A1C00162D2A377E93C860059BD59A0B8984070001556C1680",
            INIT_RAM_3C => X"A69192099BFC45A16C1048DE84217C3CAE44488081FE564ADA0852C9A4044830",
            INIT_RAM_3D => X"6FF9EA786CD6B55B4FFF2FF711898818081087294400FD71043C0428B50440F8",
            INIT_RAM_3E => X"8D00808030620AC00E4436A3809038012CB0C98D890FE01092632CC657187095",
            INIT_RAM_3F => X"A82DF593FFED92D9B7DFFFB5FFEDBEDAFC3F3B086360C056E57EB921D043C481"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1850069A48044194430C305485B37BEF1151D13C94FCC596F803FEBAE8EB2444",
            INIT_RAM_01 => X"B01360CD0188519A4CD26335919412102C49926820039D5F07515041A5246CC3",
            INIT_RAM_02 => X"ACC54067631162091E53AA03040050015A4586A11C08886904C868A288475319",
            INIT_RAM_03 => X"38D55A2A2C46394A82570C18C684FC86F0CC40F0510551154040053A39008D84",
            INIT_RAM_04 => X"55884428409359715B011009628A22818E186C68E70907043C8003D20A740844",
            INIT_RAM_05 => X"CF45EA34E338DE4239F60B133A184D8623C853604050271208510ACF50360A95",
            INIT_RAM_06 => X"B8673A802ECC50181985C86B05D744FDCB0150449534EB592ED529474452E711",
            INIT_RAM_07 => X"7788CD0715AD79822895AEDB606A5D030CDB3B5B717FC5048393DAFA3090AE91",
            INIT_RAM_08 => X"5CB6DF26BAB924D0A2571176717DB64D0CC6AAA894160F5556AA4049B722F9D3",
            INIT_RAM_09 => X"EC130048AB5181634F6D9A5400000012181803783819D3A2B064D68655050191",
            INIT_RAM_0A => X"531EF973098114D06AD6751052D1D8AC463020144003811510400FB01C0D226C",
            INIT_RAM_0B => X"81E047C1919E26F483191B40C9411B4042AB5983D1100D7E878785900D41CA6D",
            INIT_RAM_0C => X"57B0828058AC6D6B1CBA55415CC5297051AB9890D8215A0111102A0AAA403C0E",
            INIT_RAM_0D => X"B3839364357114D11A989E288902BA035B718C663F1250F08DE6152010311468",
            INIT_RAM_0E => X"7FED4489CE2A322352776E32EF8282588B6DB4EC263249364327F499A2551744",
            INIT_RAM_0F => X"6A0851B839F97D727B6C43D0F020006E61450E6147883428A0900208C89F8624",
            INIT_RAM_10 => X"4104501320B09012C410C01470224043BE1C28AC1E3063A5400A4F1D710C46A1",
            INIT_RAM_11 => X"424CF24499B5EC3246C0080A84E441D6DB58C05A551D01100F2A9049E78D1BA9",
            INIT_RAM_12 => X"A2706A5122305501044BAA80575DE9AF19190020C88106817690188022BB646A",
            INIT_RAM_13 => X"9B0F4072F6D373321C01A1A6681010804237701F84D681A9436100A032A8492C",
            INIT_RAM_14 => X"03E1CA0000060110C81029120AC050000001F8CBBBBA5BC56E9AB5B4ACD5916E",
            INIT_RAM_15 => X"010280880880CC4200A2001849A346600402868440142000320A020C82180401",
            INIT_RAM_16 => X"7853802450201C41CCC2803003A1D0EEE3A44902040C1BA48ED6A2A092A34280",
            INIT_RAM_17 => X"243C32803118120301540C058330830084E13E790181F058D19C86A01E817C20",
            INIT_RAM_18 => X"008E0000464008102043C4140980039006D0735B9466B2A8202240A24C04800C",
            INIT_RAM_19 => X"23C61A00001C466C06C000039640000180044186186186000087080034820820",
            INIT_RAM_1A => X"8009033BDCC1704E0D08CD118C6001940411555AE9F18C63140CE69D92265EB9",
            INIT_RAM_1B => X"2010C842006A030088421002910013CFE7E28A28A455542D905104D102E35917",
            INIT_RAM_1C => X"EB420140681845004AC675E1C5C203C10308001800A003C84C4E473040B06148",
            INIT_RAM_1D => X"81A0C1E09F681585F7FD9C77E0DDC8B77E791682A15A2B15EB1003BBB00DC0C0",
            INIT_RAM_1E => X"A67BE94FAD5CE6C20BC1F27E1FF988942870F0074BE069BCEF1B56A91A4B5CEB",
            INIT_RAM_1F => X"304D60417BB3518F0C0BD8F7898F542E449DFFFFFFFE3D0D1FE3E1C149C012B8",
            INIT_RAM_20 => X"634A080800041C70C8420801030D2038118600C081C56703654C80608B19A198",
            INIT_RAM_21 => X"F616808005964928884F0DCC638E230C889509A3740EDB9B6EED0C4112394F86",
            INIT_RAM_22 => X"3B5C05CE7E68182090E270C38646A4393B48741E0321AB034220056433C5989A",
            INIT_RAM_23 => X"9B224686030124C9C8DCDD88C102C928701E7CE6B15DCA3454C1183D63211D44",
            INIT_RAM_24 => X"56F7D0110788527CC8A7A08BB3F040179E1201100934289C3AB4C2A9150236B4",
            INIT_RAM_25 => X"E2698448354301C09611FE99229F43CAC27A002EACB3D6BADE76D3BE28020148",
            INIT_RAM_26 => X"1C5A473368311427011FE2108482449733CC041624040103003EA22C50129102",
            INIT_RAM_27 => X"804062991CFF9E83283F2C31124C0824208C49261841924466234C803E408D80",
            INIT_RAM_28 => X"78B6DBC3F054F02078201E08F010C2C52F96058665311141C004A4E08C492610",
            INIT_RAM_29 => X"06C55B5412224DE8D92E89AD5E8CDB6CC9D51A8B6D0984AC971AD56A6E0B445B",
            INIT_RAM_2A => X"770F22127AFB1C37324D6EB98CAD86BFE18120499892501892AC34010C9C4548",
            INIT_RAM_2B => X"0B97F7DCAA0041FA05CF7BEE5500201DD54E7A7AD7198B5C919A6CA8C1CC6272",
            INIT_RAM_2C => X"AAAAA5800204840001B4F7BDF62B8999FF64F714DBDDCB3A173DD60ECDE98074",
            INIT_RAM_2D => X"FDEEA6420DA65C2B7179A9A7FFD42BDF90816B4F5AD6886B936F78C90862DAAA",
            INIT_RAM_2E => X"D60894555922E462034B5AAD5EAB57AC8100D686B4E33254230FF3F5B42D9B74",
            INIT_RAM_2F => X"D4F7FD662E0F16ED4604750A9052D6CA390302180C5BC9515396405553960053",
            INIT_RAM_30 => X"600E926835238221F4A40090029B95F26233A94C1FBE261BD3732D91332F5CFF",
            INIT_RAM_31 => X"D33623811F86346DCDAE0F800007AC7DD831824C453E68C0939DD795744C59FB",
            INIT_RAM_32 => X"DC560C79200A6820032707125A40638C5A3206259222218F16F04F312488B86A",
            INIT_RAM_33 => X"A20E19B4214971DD6EA964205A2127180319CCE994C4C9362C44A719A668AD92",
            INIT_RAM_34 => X"481F88B43292D09500A490842B26239A92224DA8856C8930C5EED1BC09B31843",
            INIT_RAM_35 => X"269244034E08191080552A5CE8289802A6061146C186EB7B44C18688AE688D98",
            INIT_RAM_36 => X"6A69881020DADB1AD00CC4800145270DE85DDB6AB2ECF68B1941344F6B1AD204",
            INIT_RAM_37 => X"0E4905360440904B00091A3B3F9464E229D69DC01808F08C1B14271D51BFB6DB",
            INIT_RAM_38 => X"F4F605E6EF0C55720044D4DF9FEAAB02B7B6A4CCB52F6A1F16405D68AB3E708A",
            INIT_RAM_39 => X"8BD2886D2EA71D13B0595AD6A56A5AA17ADC69A7BE1CEFC5B3FF74F1E86745FC",
            INIT_RAM_3A => X"B42825EA097B71315B5CC050C3143243240B12230A46915C0EAC07595223198B",
            INIT_RAM_3B => X"9C7428E124F409014F73112F6E223E2832E44AE3C53B2A33CA2F3BBB510DB6EA",
            INIT_RAM_3C => X"F490927912AA10C6914749DFC53B0180327741F900070C75124259002464C310",
            INIT_RAM_3D => X"51EB5AD62637ADBB4FFFEFFBA34FA74B4E180F81164D4954046A1210830C10F0",
            INIT_RAM_3E => X"0929A90CD16A46F1FE4EC4AB2F50F9932CB0A90C890FFFB892412482024B332A",
            INIT_RAM_3F => X"EA0B2DB6CB6492DBF6FFFFB6DB7FF6DEFD7F795C51627F14E92419320C60A484"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C44AA1259758B4690471C4C833E0FF7DEAAB8429FDEC44155B12051142451205",
            INIT_RAM_01 => X"03E407125A0422009004082040228445C0A26607D5E43E10B82623220B899134",
            INIT_RAM_02 => X"9022880010E48790015052C03AB08580E01A2B4C01033194ED71959104000006",
            INIT_RAM_03 => X"E357EF662CC6610AD06A4890851084101100B000401115445151110944805210",
            INIT_RAM_04 => X"11425832C48450401D0018A1009ACA80C228A40B0440A204204658654DA19624",
            INIT_RAM_05 => X"EC59B327446ED919B9102E6664C337242015C288608105A348004B6C05254A31",
            INIT_RAM_06 => X"21041059B320E153421229045514542C295405544000448DF32E93F1E402A79D",
            INIT_RAM_07 => X"2266602135B583C72914000A048A500008010909610410231B7B2854EC0CB37E",
            INIT_RAM_08 => X"58924050482D045A04D6D540010492420960AAA9358081554AAEC010210B0704",
            INIT_RAM_09 => X"455140646188436DA100A0894C554501710740810262300AC22112708E000093",
            INIT_RAM_0A => X"1ACB3D40607113426C5D8CC74014439039CE6A0D1590020A0C9E4C44380D3141",
            INIT_RAM_0B => X"0C836124CC910292224148CE000148CB22A902985133C84830180E09341210B3",
            INIT_RAM_0C => X"D22650302C24359C6049540141140C9484A2120846C54836900CAA00A0810802",
            INIT_RAM_0D => X"001202C99A24200CEA0080299594A82C54139CE39F1A007000A840444D883081",
            INIT_RAM_0E => X"00241B26846EC90949998850183B2800000002008A00003200200211D395307B",
            INIT_RAM_0F => X"6000C082AD44830001248840D99800684272B088890890CED42004002014484E",
            INIT_RAM_10 => X"E2340464A2000ECC93DA394007204358B4C0655A222112080040230046B00003",
            INIT_RAM_11 => X"4208C0300801BD0C2048182A240010DB6D8C610A544D51473044605203264AF0",
            INIT_RAM_12 => X"700A0C98B2B75E68A198BB0A998090304383840D1C36485997788CE628201188",
            INIT_RAM_13 => X"40401A11124014848522929364014AC886C42D240518C02930084248211D1471",
            INIT_RAM_14 => X"6B042100888A4A46A346894C45410000D41918044444481400025296311A0800",
            INIT_RAM_15 => X"21A800B9CED912B5BCE60400B6A54888119AA2BC8C011C6022A02AB04C85533C",
            INIT_RAM_16 => X"8230411330135336111180026AFA201111491256CA5A4000115192AA82982C00",
            INIT_RAM_17 => X"C66582A919320603155988CC148460124054810499790CC9114BC922112B0B7C",
            INIT_RAM_18 => X"8021100026444891226A886663424101A505667A004494C30CA08C4923324A0D",
            INIT_RAM_19 => X"4088B3C0D695E35C05155578288AAB22022235441041042004424E0118000002",
            INIT_RAM_1A => X"004C19D3618064374E010002108406C00000001C23318C6340068C8C902354A9",
            INIT_RAM_1B => X"04848210806049210084210300002A20124000000A8023D202086059826E6815",
            INIT_RAM_1C => X"1D8001800059018000CC2110A6911A22C58288A200C40080081826E762CA6594",
            INIT_RAM_1D => X"508921880B4C158831FEAE54D825003226A93313A3D9EB35289A14444D626911",
            INIT_RAM_1E => X"846C4108A2C138E6410986710012DD1C3870F0269316A889131A7668BABF554A",
            INIT_RAM_1F => X"11A940F1DAB0FFE5084490238B82260C9CA8000000021E1C0FC3C3C1D9400234",
            INIT_RAM_20 => X"A583040000042810008410819E11642944D4A9A395094A530146D59541C93212",
            INIT_RAM_21 => X"C02601100184C11892011224A6C40976B3C0200F008000200000D9C718D0EC28",
            INIT_RAM_22 => X"0B140508480A084804401940D524460C1240240C110180031000000CB03482B0",
            INIT_RAM_23 => X"92282366080A4A14616A3099C125902A20229DD76B397B7D9960402948321046",
            INIT_RAM_24 => X"425246286217621C940901504006232000084B08F120280410864400232AB436",
            INIT_RAM_25 => X"1CC93320027409CC36266C8803082C5C2D17AA32BB84E000000004004050A508",
            INIT_RAM_26 => X"852CF199BE834159D49826484C202246682124911821646ABB8548CD652064E9",
            INIT_RAM_27 => X"193BB92249A802E49687C214C93830C99C6336D8408364C84C9891350914264C",
            INIT_RAM_28 => X"228003FBF41962698B0262C015102F0C8000180103E064326BB90C2C6336D841",
            INIT_RAM_29 => X"207310006DD000482C7B449185424000A00B0F4000A8A2663D8918D904613309",
            INIT_RAM_2A => X"8CE2F48C061C808089B7209441A4000101088030800C07822448A2A6E801B104",
            INIT_RAM_2B => X"0BB3EC230B08CA1696DA44139796770A802730858DA4604834060030042118CC",
            INIT_RAM_2C => X"CCCC780000020C0001F5F7BB09CBCBBBFE0948A106B226485775E267DDDA7C2D",
            INIT_RAM_2D => X"9420B01ACE029D2534F80E1249432540090DB9006318408D4861326C205800CC",
            INIT_RAM_2E => X"31002683224B99313181C8844A25108C0C13721B901300213C248A50C0220C12",
            INIT_RAM_2F => X"198A0D06C19B739618318C70089A0812E41975A4B46605A2CE71B308CE70C34E",
            INIT_RAM_30 => X"0D49B0647240245814A030DB21089408D9D93A550AE3A8CC931A57244D0388D0",
            INIT_RAM_31 => X"82899900622890A49448D2000019BC2556DA2911131089719CD3B00812828030",
            INIT_RAM_32 => X"DDD11304D7449208C18211A9C65D3894C0CF06F2368C9C103024AEB78DA33064",
            INIT_RAM_33 => X"B1A0CA851DC9A000033620A5009DB0E73998C4EB2599191064C42319B7A42492",
            INIT_RAM_34 => X"99520042C842168966F3344838DA6DA9A6DD64992C0308876220D80D088DA9B8",
            INIT_RAM_35 => X"A3CCC8441261CD8D2E87024C01040A010F89E5F952B44CF2D214E06116946245",
            INIT_RAM_36 => X"00434810294E496E40108088849730640A10001B8CA410B9392313E0220A14D9",
            INIT_RAM_37 => X"800012C40E16256229244D82401130AE22223081CD90D990C89565A231000000",
            INIT_RAM_38 => X"934A1251839C85D5FD6D61A880604302131982C0DC2538339C44A1CD2E275A50",
            INIT_RAM_39 => X"2259B240F90FF0D85819C44A971CCB990E30228A11B180DC8D2521449B304D33",
            INIT_RAM_3A => X"566AF566BD5B115400023F160C4509844965CD11509B935B693C442D5A42AC08",
            INIT_RAM_3B => X"0005AA1D9005BB6450CD9D3032003666B4211AAD4C482910409801CA3700D251",
            INIT_RAM_3C => X"76D307782002036257E9D8D29AD45668CA1CC60475582000664E354ED6222DC8",
            INIT_RAM_3D => X"55212C410012846909242490C001228498B204516648AAEBFBA966B5835864D0",
            INIT_RAM_3E => X"D633333BC060331008032656E9532225249029BD8319242800100020AA10492A",
            INIT_RAM_3F => X"AAC01801A6C00092D20082506816DB4C1224303792CC68719009914E56B948FA"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000200002CFB7BEFFBBFAFFEECAEEFAABFEFBEAFBAFEB00E",
            INIT_RAM_01 => X"040808200440044022010042044108020000000000001C0F0010100000000008",
            INIT_RAM_02 => X"0110010088001002002400140008005001200002002402020002020040800840",
            INIT_RAM_03 => X"F600C104D89DDEE5D59442008460FE002012060BABEBEBFAFEFEBE0000280028",
            INIT_RAM_04 => X"264FB3E5A357BF7D64DDCA53FDCBEEB9ADFABBFEAEDB46DEF0B60BFBF88A8ADE",
            INIT_RAM_05 => X"D4F51120C07ED391D99062292D63AF0473333095951E7965D57CF60CD7A4BC06",
            INIT_RAM_06 => X"24AEF4D4155EA21839D92EFA4DF7A487C6D57D7F9B3CB95A55204208B0FEE51A",
            INIT_RAM_07 => X"AB30FBB396B5A0D3699FC93FD64FFCADBBB7ED9D97BA8BC6BD752CF560CA158A",
            INIT_RAM_08 => X"65B6DCCD453B3CA5F67CBBEFDD96DBECF0D5AFAF1A4C6F5F4FF8F81DFBEE2364",
            INIT_RAM_09 => X"DBFED4C7272637D25E93F0B9A0A838ECA49E0FDDE9022ECBE9FD1DE99E0A23F9",
            INIT_RAM_0A => X"9E1B6FD51A8B84FED5ADCA677F68FB758842D07F4BF77B616582DDC0F3FBC1F5",
            INIT_RAM_0B => X"A3AC8775EBD7FFF946B69FB1A8569FACBEBEEE56539ABEF7AEF0BEBF6F98C44A",
            INIT_RAM_0C => X"1CF1570AC1BE35BC959F74A1F1975F2FA1F19B08D1975E8E38E33A50F0A03577",
            INIT_RAM_0D => X"7D79EBC33CE640443B1BD168F3D5D7BA6AD18C629EB7AC7DC919685500421004",
            INIT_RAM_0E => X"FFDF8B14BDF92D43E4CCD05FCB172C4FAB6DB44ADF6DB6E97BBCCF55180D1C0C",
            INIT_RAM_0F => X"F0C3E3E118FF0E8DF7DF2E6FDC073559AC0D63BA3DF185012CEAD5FF9EFDB944",
            INIT_RAM_10 => X"0F1978C323801120CBB39460C6B06E77F6B57EC387BC5FAFF57076BDDB609C4F",
            INIT_RAM_11 => X"3188F27922432BE1BDAFFC101A980D2000110B45E0107C7E040C05E93E8194C2",
            INIT_RAM_12 => X"0B6A4526C5ED107DAA85143AA01D4540C0202CDBA16CB9A6A92205F28F3278CC",
            INIT_RAM_13 => X"E4F8143F3B64BFED1FFE6DF7E343FFFEB87B877A28CA6B10AB02160BDD55B400",
            INIT_RAM_14 => X"7F09C152667936FF03D3B468477541EAE1EBF5B11112DB164D2652DD610A8A4D",
            INIT_RAM_15 => X"96443E04270B77ADFDC1F2D3911C39BB508D443EC75E3D4A58F06BC8FD7D5104",
            INIT_RAM_16 => X"9CFA7A2006B96191F7356BEF2D963AF7375FF7AFF936DB6B782C4F0F1C525C6F",
            INIT_RAM_17 => X"9BCFEEBE7DC6D2ED75F8ABBF5CDD6E3F59093E7FF56A0FBD9DC979596FD78507",
            INIT_RAM_18 => X"74D35DDD98D64C993266EF9F3B498B5C7DF9E2D7755DDBD14EB4F17C4D7930FA",
            INIT_RAM_19 => X"B2F83EC0D6BC68440A55541EFA62233E79999D75D75D75FFF7267DFF3AFBEFBE",
            INIT_RAM_1A => X"45FF3A776DBDE24933FB4756B5ADA87FF7DF7DE2212F7BDEF54F85FFFF76FDDF",
            INIT_RAM_1B => X"BD6BB5AD6D5556EB45AD6B6A5DDDE660062FBEFBF3FF36E9596596FFEEDECF3F",
            INIT_RAM_1C => X"882F550EE5D7BDEA7EA5ADCFBE8FFB162C476DB6D69553B66F5FBEBD7E96DD2D",
            INIT_RAM_1D => X"5587A967B2DB5F7DDEB63E88CF83BAFEA7FE8B5E3B3C468B1A63C66661C70C98",
            INIT_RAM_1E => X"203DF04769B9B8FA6B19305D81B051D7AF5EAD64D27881BD14B68F8E37C6F9FF",
            INIT_RAM_1F => X"9C7FE033C717B56F6B71FD79D1569D5C7FDBFFFFFFFE3C3C07C1E2E1C04150A4",
            INIT_RAM_20 => X"9316CDCD7D7FDFBD75ADB5B5EF9D5A5F417FEC3BB596F6D7E6EFB32BD3D36874",
            INIT_RAM_21 => X"CD6F1B6DABDC56DB77BAFE0797F9E98F55BED1B6FF620019244BFAFB6FD7DDA5",
            INIT_RAM_22 => X"134A061088B59EBD78D9FCFFE4BD1DFB36DFEFFDFEDBD6B7854B6A8B7B27F8E5",
            INIT_RAM_23 => X"5242465D0F0D034082FF37CE7FDD115C681E18DEED0A5BD5B8DF0DFBE0F8E1AB",
            INIT_RAM_24 => X"80648D05C71DD02606C747E004FD07803FE0104160ADDD4BF7FFBF7F9C6AAEAC",
            INIT_RAM_25 => X"18B943D12AF03609A6BC5F11DE4D8B97F86550674E631610421011840FAF06F5",
            INIT_RAM_26 => X"1E68A640C138B9398BE7C5F48A29C12B07C6AAAA215110131543011AA8044244",
            INIT_RAM_27 => X"0096260424BD77833878187803838011489C260B8FA888B2E245020A2023C183",
            INIT_RAM_28 => X"30DB6C0002318D57326CCC8BB80389E3494D435C3A010BC1D3420B989C260BBF",
            INIT_RAM_29 => X"C0A7C3DFCB3FC195C01D1BFADD1F2DB703E2A9BB6D5063980EBFADD7CE4671B2",
            INIT_RAM_2A => X"1CA7AA9D307088008994091DCFC810BE68A248AB448F8A91189F859C171F0EFF",
            INIT_RAM_2B => X"6687402424242402334D721212121201D5AF7A0C029C018CA4A7044218413480",
            INIT_RAM_2C => X"5A5A02000000080001B4929900000080FEC0F08430C8010A850EBFFFB7B3B004",
            INIT_RAM_2D => X"E80DC686B7EFFA466815B7C49084809FB4EB2066DFF73BFDF6C061598BC5E85A",
            INIT_RAM_2E => X"A7CCFDF8FFF638B56F35031184C06333A3EB40F2064EB7E5CF893421BDA4B8BD",
            INIT_RAM_2F => X"B4344E2FA7FAC42B7BAE383B9EF47FBD8E56C3F50AD09ADD1CA5BEF71CE52C9C",
            INIT_RAM_30 => X"6BF3FFC22088018298C3C924CC81F5B0595D6BCDEEF2D9EEB4772B12322B1540",
            INIT_RAM_31 => X"A0C9CD6ACC920A08C192BA4554317AEAAF9E103088F6CF766ABB884000200033",
            INIT_RAM_32 => X"0AA7720088FC4C7123754D28E59B05CE778BD8221D8D82B29DE80C410F6372AA",
            INIT_RAM_33 => X"75E63EEE3FF4F0008BBE022C2110E24288AD56370B8B0E275EA8E738E090C9A6",
            INIT_RAM_34 => X"8E3E991546B7BDBFF332188C091BDD7F7DCADFF51A6BD9B6578DB5BB59B96F29",
            INIT_RAM_35 => X"ECC86C4759574BAFD7E8FD8FA830F0126BA8EB7971B3D8E40A3CAF1CED59563B",
            INIT_RAM_36 => X"6E51355FF08891B81A8777E66CECD31FDC5D9B74917F7DDFD769EEDDDEBFBDB0",
            INIT_RAM_37 => X"FA79FC2CBD696196B6B06F5E498C38F10838867F0BBF9441D3775F678B4DB6DB",
            INIT_RAM_38 => X"2515BBFB3F4765FD5F5F44B3E05F8CF847302DAF814263067F91777BD7E2F5BF",
            INIT_RAM_39 => X"1163511C32FB622ED76794810C5816263C86C10424260EB022423E993E61BE63",
            INIT_RAM_3A => X"556EBD7FAF5F737530083C29F0FA21D0990A08337DFAF96341FAD0BBF7599AF8",
            INIT_RAM_3B => X"B5EF6CD36DEFFFFE86C5AFE3E2E67532CA510EEF69555131F2A6C38A9B82A42C",
            INIT_RAM_3C => X"ADBC139F9FFF2757FD6AB7A3A034845132A154D8361AB00063F3BB5D6DEDD835",
            INIT_RAM_3D => X"D5821C8D666308001000401ED843CD18481268D3C405FFFAEAAFC01141F8C056",
            INIT_RAM_3E => X"C86260436AFD427DF0EA555C77BDF3DBE53EDF4FC972301C0248049104C221EA",
            INIT_RAM_3F => X"B82491B7348DB649D249B49A6D3492688048624C698A60C42E1C2105AA422439"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FFFFFFFFFFFFFFFFFFFDFFFFCB2DB25B01052BD644517A1110FC410100044FFE",
            INIT_RAM_01 => X"FBF7F7DFFBBFFBBFDDFEFFBDDBBEF7FDFFFFFFFFFFFFE3F0FFEFEFFFFFFFFFF7",
            INIT_RAM_02 => X"FEEFFEFF77FFEFFDFFDBFFEBFFF7FFAFFEDFFFFDFFDBFDFDFFFDFDFFBF7FF7BF",
            INIT_RAM_03 => X"17FD6A32664A570E00E44C98419478F81F0CF86001540155005540FFFFD7FFD7",
            INIT_RAM_04 => X"30405D781130C6602D1011012682CA918024C04AD5048300009146DB0B445188",
            INIT_RAM_05 => X"42DD77038752970B90F0211454D17B8022C970B0C0500B9100010A4800240291",
            INIT_RAM_06 => X"31550A156AA1C0121A92A82D4D962055400000064020820EA2261266D406B404",
            INIT_RAM_07 => X"1008A52396295A8E01B426C004A80300AA01125B8118900340D0BA68F8D6AA33",
            INIT_RAM_08 => X"60B4992050AF34C002582202214936414D4100A0A0D606000CA46D01050BCE97",
            INIT_RAM_09 => X"01685428DAF5A00284488A0D20802080480C07A93BAAC322432150F7BC000039",
            INIT_RAM_0A => X"185E4CE804210300281AB9DD40A04208D6B42A2554A1D0C8C31186B01EA0B725",
            INIT_RAM_0B => X"48C6218488900202C30A0814100208094680011084309A00215B438030538434",
            INIT_RAM_0C => X"E92460853D25697A282955554D54845211A00288540549249088AAAAAA140298",
            INIT_RAM_0D => X"A223232B33155E9112808A3D8940002D42308000910954008D0445044FBDE3FB",
            INIT_RAM_0E => X"000445A9E70456234BBBAA601C81880EBB6DB4E0EE3B6D8452113088A3C7B0F8",
            INIT_RAM_0F => X"2186008A9494E45B2104291A31DF156603B8095016889077042550F60CC7846E",
            INIT_RAM_10 => X"F2AD0035120A0C5496120040102847408C842F813EA81CA1550C1915500A3118",
            INIT_RAM_11 => X"21441B46D1207403100B401A968D4956DB4AD01A15150507B97F7A82F59F98FC",
            INIT_RAM_12 => X"3B3A0B97231FFC6C01CCAF4A5359502E59594400FC0604175ABCF855A02251AA",
            INIT_RAM_13 => X"5B234010D6DB508004110333194084009F08850004108CB5906522DB0C954B35",
            INIT_RAM_14 => X"05D9C150444450522B52B45D56D5406A5549681BBBBA5A5568DAB5B2A6CD5168",
            INIT_RAM_15 => X"82AA828D31448A421A77105064B364400556A2B0AA011A500A0A0038003000A2",
            INIT_RAM_16 => X"7C510822AC282AAA88C0828505C0A0AAE0A1405244345A06C6DAB0A09AE92EA0",
            INIT_RAM_17 => X"311486A829081205154D0EE01320440088B5AF544798BA09551F26082A29521A",
            INIT_RAM_18 => X"F46B555570224489122F4F5065C343D43B553401D77061EC24A25022481490A0",
            INIT_RAM_19 => X"51E622804200287C0BD55408F24001013BBBBDD75D75D77FFF27B55526EBAEBA",
            INIT_RAM_1A => X"01F51241BCED36403368457084200F6AA61861804A54A5294000282545890024",
            INIT_RAM_1B => X"AC42A108400A496844210801C44410A039AEBAEB9555004873CF3C4E2C0C1104",
            INIT_RAM_1C => X"4B0554CA0D406C2B2607150971C9CEB972E0F668077550E2210931D576F40DE8",
            INIT_RAM_1D => X"142C690405214088D6819618650CEB844A5594CBD3E86D76F052D555513AC959",
            INIT_RAM_1E => X"00198080C0C574A551A947535EB888C68D1A28251290A90C45017AF428050500",
            INIT_RAM_1F => X"A0E00027DE1696A06E63409482891226D800000000041C3F0FC1E3C2C0410024",
            INIT_RAM_20 => X"44C14545555281003C608C0190259F255150AD6A544B09546310556A8AD090C2",
            INIT_RAM_21 => X"B13489B4810F6A4D180412AC44924B2412C0601301A200100236576DB4FB6B22",
            INIT_RAM_22 => X"1302054AB2588058B02F40AA061232A5080A82AA00492892162920212074BA8C",
            INIT_RAM_23 => X"120222D0000000857B968EDF52674128300372CFBDFE4B58A4AA1E80038194CC",
            INIT_RAM_24 => X"C2524EB1C387F02E0445A01FF802F87FC001EFBEA8C0893149081402A8002020",
            INIT_RAM_25 => X"7EB51648137152BFA42FD000F2DB6A8A6B22AA2E2B71400A0000010A04D6A218",
            INIT_RAM_26 => X"8DFE52B17AF0DD0E773576906C35265A796228A10F396028A9A83A791502E5AB",
            INIT_RAM_27 => X"DD695AAD19EFAEE1FBC8B6366A572CB5A847E59649E25AD60C6357951575ABCD",
            INIT_RAM_28 => X"2FA490000235E75BD387F4E17551EACBBF8B96CB22585710AD96CD7847ACB259",
            INIT_RAM_29 => X"60569004C88300F8782A09AD190E9249F8C28AD249B8A2DC151AD18771693549",
            INIT_RAM_2A => X"2F8260EA3E2E7C00A34F649543E4A06B200C8421180A590E876DA2ACA487234C",
            INIT_RAM_2B => X"0918BFDBDBD9D80284828DEDEDECEC01DDED602F180CA8CAA0C3028404A50AA2",
            INIT_RAM_2C => X"936C73800000000001B4929900000080FEA05A016CA2A4581231400000000005",
            INIT_RAM_2D => X"1424C7541D24DC6531301D124843614F91823B025294094F92612AE95C82056C",
            INIT_RAM_2E => X"712224807B6A9D4175E5D984CA61329489367633B03652510A249210A43D8E24",
            INIT_RAM_2F => X"7D827924D89753829702C454091A1E9AA513652E2D7629EACE31643A4E30804E",
            INIT_RAM_30 => X"2919303DDE77FC7D5FF036DB337C34A6263BAB45B983B4DDDA1827870C4144EA",
            INIT_RAM_31 => X"D0ABABA05F96A62484B0978D103F287CD6A5A96D525EAAF929D2033EFF9FBFA8",
            INIT_RAM_32 => X"90ABAE002246949271ADDA5B9499611811FB8846A4ACB0DF0407F3C2292B280D",
            INIT_RAM_33 => X"812E1220191007800CC331173998335B1BA1108789D952061C20442176404924",
            INIT_RAM_34 => X"5C152244B098862864B6A00690766BA9A6A86A98ED07888FE4009009088FA1F7",
            INIT_RAM_35 => X"0ADA8620164BBC09048040C941C73A8B6BAAD9F5D091EED1D6E5B6C544944589",
            INIT_RAM_36 => X"0563981031CEC80EC00C442AA794570940184019036944037A33B06E621084D5",
            INIT_RAM_37 => X"9441015B5632D56F93275BB15781F46006D69271BC12F006E9356B8E21A00000",
            INIT_RAM_38 => X"91C01EE59D1665DDFFEF74519F40A602129D8494EC2538539C842DCD065B1010",
            INIT_RAM_39 => X"A8C99E07F86B5809B8314240851E42812250E082123395DD89212C449194C953",
            INIT_RAM_3A => X"FE7AB5EBAD791915E8429DF445310A45B53255115895D963E728402950488C6B",
            INIT_RAM_3B => X"06A180F9A6A1B365822209383B48ACFACDE90A2BC4380910909268983BC3F28E",
            INIT_RAM_3C => X"F4D2175AAD1102C63500DAD2D0938500E20F4153140C28005F46206C66344E90",
            INIT_RAM_3D => X"81E50F41005084C909242497F80111FEADDD04007000EEBFBAFEC1022907F4C0",
            INIT_RAM_3E => X"82F0A017584A1793582ED80536903849AC90C93D0B292A9C0008001100C10A40",
            INIT_RAM_3F => X"FFEDB493FFA49249F6DBFFB6DBEDB7DEB024382721A815D18513681E86168452"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"22411114482102912242088926DB4924ABFAAEBFB8BABEEEEBAAABEAFBFEA00B",
            INIT_RAM_01 => X"400080020000800200100800144108922449249249249E9F8911512422491108",
            INIT_RAM_02 => X"8000100800100080020002001000800040020200020040000410001000008000",
            INIT_RAM_03 => X"43AAF55552A97AD52C714A94A55CFE000000000EABFFFEAAAAFFFF8820002000",
            INIT_RAM_04 => X"8ACC9D7A9436AACA86AAAAC64D17E160DCDCD9B260599735B4255555CAA9552D",
            INIT_RAM_05 => X"DEBDF72E9552DE8FF1ED555750557B8551A3B2B16AC567B552AE92AEAAB6B9AA",
            INIT_RAM_06 => X"6560B9555DE8AABA2707A24F532C8AAE962AAAAE5C8A16DCDDAB5AAEAAA9D71F",
            INIT_RAM_07 => X"AB2BBB00A95AE25555AB193260E37C5F41DB648453265D9F97D7BDA8F86D5DAB",
            INIT_RAM_08 => X"8C4924897E7CAAAC56A2AAA4D83249CE916455562AE8F8AAAD54E2D55B6366E0",
            INIT_RAM_09 => X"C8BA2AAE758B5740E313B5D02A208A00EAAEA9B062FBB6C8E2EDC6F7BAAAAA4A",
            INIT_RAM_0A => X"384B5C5108AB979368CAAB751322CBB62D6AE558AB162AAAAAD558C5395DB6ED",
            INIT_RAM_0B => X"8BA6A764CB9BA672973A39C5895639C171566C562AB8AA24ACDB8FBDB983D697",
            INIT_RAM_0C => X"04F5560ACF8CDAD6BC990AAAB1519DB6D454AAAAB000BA28B980855555CAAD64",
            INIT_RAM_0D => X"519E86888AE0A815705D945563901A0D19C94A52963A2A79207172E540000000",
            INIT_RAM_0E => X"A4ED9F3E9CE57DA8ABEFB91BDE3321414492491CAB04926295ECCC77DFAAAA2C",
            INIT_RAM_0F => X"6451CAF07BED9B24DB6CE2659954AAE9F2AB36EA09156E7562AAAE3BBAAC310A",
            INIT_RAM_10 => X"AAAAAAE508D47D55D798B10AC6050B1BA68D7D50BF75555CAAE5662A0BB00C07",
            INIT_RAM_11 => X"5288E4B12A4399EE8EC0B865A812D42DB6D5AAB5CB42AAAEAC5F556A8CAFC55A",
            INIT_RAM_12 => X"54D556AB554EBB5558D353558EC4015EB8B8AACDB576B138E1AAB5555544B3A2",
            INIT_RAM_13 => X"C4ECB9B73124B7B67DB44F7726AAB54CADE64876AAAD534A62E315D47310E45D",
            INIT_RAM_14 => X"5103D6AAAAB1572CAAB54A5D55EAAA95CAAB99C66664A51096256A4E69BBAA96",
            INIT_RAM_15 => X"A85555555555DAC63ED55502EC468CEAB155557CAAAABE5555555573C94AAAAB",
            INIT_RAM_16 => X"C2A2E2AAA94A82AA5D95957150EB355D976CBB2C9142A5B131AD6E5545161C4A",
            INIT_RAM_17 => X"ECEDB1555832B550AAB9C1DD84D572BB654A50ADBB6A6CD943C94DAA85962D6C",
            INIT_RAM_18 => X"0AE8AAAAAAC54A952A522A861DAAA92AABAAE73A28CE9AC15C85C5EC9571255D",
            INIT_RAM_19 => X"EE5832234A4A92A013800516F0AAAAAC4AAAAB2CB2CB2C800552D40011145145",
            INIT_RAM_1A => X"02D8B8726092E5804295B28B5AD5568008A28A2733A318C62AAECEF89F3E7CF9",
            INIT_RAM_1B => X"52B41AD6AAC55495B2D6B5572AAAC710365555557580245A2AAAAAFB94C74CBF",
            INIT_RAM_1C => X"5AAAAB95D2B9D39099C6E3C32C9555AB56B2B0FAA8CAAA9D585CACE669EAC3D5",
            INIT_RAM_1D => X"5D8AD5A0B346ABB431AC508080AB1462244C830773B854C112081575742AA155",
            INIT_RAM_1E => X"A64D994B48AD76DD5D55D566BE1389B162C587575BA8D53940BA6EDC33C67BCF",
            INIT_RAM_1F => X"9119E10F004E20029954D1739B170E5CAED9FFFFFFFC3C0E2FC3E3F3F84252B4",
            INIT_RAM_20 => X"179F3AAAAAACF9F9F2D55AAB92102D58B42C55D5CB16472B167E8B5552E3B3B1",
            INIT_RAM_21 => X"CF2659248B9DE61D24D26B2B16C9AAA655CAE52F2B844901244BD9E79E99ECAD",
            INIT_RAM_22 => X"AF230339C8B95CB962E9F84FCC8C0CF8BA47E4FCBB499793555922DD33318234",
            INIT_RAM_23 => X"5B5556BD5F5F274A9596AD57F34988D1705DC520C0D41DCF184F74D9EE7072BC",
            INIT_RAM_24 => X"52D6D7BC6F2FF2F8DFAB9000000000000008000029AFD7C9B9699B14AB557171",
            INIT_RAM_25 => X"7E7E5E4D7BB7F07F9297FDDD9B4D3A0EEB83FF6E7F74773F5AD6D7B76E7CF4AD",
            INIT_RAM_26 => X"D9EE78FDEBF2F16AFF82B7D1CF3873537EB62EBBAFB07628FFD57F7D9FB7F5FF",
            INIT_RAM_27 => X"5D7D5F2E5549B4F5FFE4BB66FF562EB9CDEFFFFE7D235CFB0CAB971FAB9F3E6E",
            INIT_RAM_28 => X"5FDB6FFE64D5EB5DC3AB70EBA7FB3BCBE9AD174DF35D561ABDD70FBDEFFFFE71",
            INIT_RAM_29 => X"B47F71FC5FF76899FE335BADFD5EADB7BBCABBEDB6FEFBDF19BADFD77FE1710B",
            INIT_RAM_2A => X"AA0862FF4E8EB634AB9769BFFDEDD695722E8EA32DBE7BBBD77CE3F7FCDD774C",
            INIT_RAM_2B => X"412D3FDBDBD9DBFE00000000000000F15FBBDAA94A3DAB5795F76FCED5AD6AAA",
            INIT_RAM_2C => X"1C7008000000040001B5929908080188FECD3A2D75ABA55ECA5A7FB7FFFBFFF7",
            INIT_RAM_2D => X"4D2E1A1845B68DAD76916792DAD7E95FD9CCBB777BDE2CE8DB2962C6A908818F",
            INIT_RAM_2E => X"13BFE689FA66B97573D9DAA55AA956A385BE76D3B77E3B65CB25BAB5B6E6DEF4",
            INIT_RAM_2F => X"DD96E974FFD2538BF316FD5FDCFAFED9AC5F7B34F8F65DFBDE13257FDE12E94E",
            INIT_RAM_30 => X"6FA9A540208801001F00000000001CBABBBBBA6F0EF7B5DDD9390F952BE74994",
            INIT_RAM_31 => X"D2ABABA2C630B8EDDD82FA72101FBCEDCC8CFD67FBB0A33DC9C3944080202032",
            INIT_RAM_32 => X"4EFD2682AAE8D5D75B80D1AAEC192B9C72FD13763C8C95D31C88001BAF2332FD",
            INIT_RAM_33 => X"B5E07AE7BF65000080000080000500C72A9CE67F2F991DBE7CEEB39CB27E8492",
            INIT_RAM_34 => X"1DDEFF7C4F9B9EDDE7F63EE3DD5369BF2689E6F1FC4F1DD7E1A5D89D9DDFBB3F",
            INIT_RAM_35 => X"F5D8E377F175FDAF1789BC5995D74FDF65AAF9FDFBD66ED6DAB466ADF45D7E79",
            INIT_RAM_36 => X"49E2E7EFCDDEDB9EDFD7776EEE8D903CCF508933DC6D5CCB7863B6E9EF3B9ED1",
            INIT_RAM_37 => X"D914637DFE72E46E3B0555EC4C1574F22ABA9177BDB198D7C99FC18213892492",
            INIT_RAM_38 => X"91C5DE20819645FF55576140C0EF88FE973C8E8EE46D6991BC0463CD163739B1",
            INIT_RAM_39 => X"ABEB1F6CF8EFFAE8D3C742D1BD5E568562972BAE9411AC9DA96B7CD4B9543D13",
            INIT_RAM_3A => X"FE7FDFBFFFFDBBBF339ABFF6C523AA45D9795DBBF193DBCBEFBCE6ADF94BDCCF",
            INIT_RAM_3B => X"3E67BFD5A6673F451AABAFB2773FF4FF9DE08A3F64395BBBC29613AABBEDF662",
            INIT_RAM_3C => X"249AC66DBBFC4663DFE6D0D5D4A42541F72BE55550BB27FFCF6F77CF6674CEF1",
            INIT_RAM_3D => X"7F2B7CD56AF5ADDB5B6D6DAEF35B1FFEB9F7BDFAF24DFABEABAA53977DA776D6",
            INIT_RAM_3E => X"9AB9EB53E8EF5738AACAFD147F99326DA6BA4D19A30B5501B6D36DA6EF1A6BBF",
            INIT_RAM_3F => X"B8249801B6C00000D249B69349B49268D4ADF32F60886A518E77737F9ED62DF7"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_basic_kernal
