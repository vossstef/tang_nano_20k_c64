--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Fri Sep 22 17:00:33 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_cart is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(12 downto 0)
    );
end Gowin_pROM_cart;

architecture Behavioral of Gowin_pROM_cart is

    signal prom_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= prom_inst_0_DO_o(1 downto 0) ;
    prom_inst_0_dout_w(29 downto 0) <= prom_inst_0_DO_o(31 downto 2) ;
    prom_inst_1_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= prom_inst_1_DO_o(1 downto 0) ;
    prom_inst_1_dout_w(29 downto 0) <= prom_inst_1_DO_o(31 downto 2) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    prom_inst_3_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= prom_inst_3_DO_o(1 downto 0) ;
    prom_inst_3_dout_w(29 downto 0) <= prom_inst_3_DO_o(31 downto 2) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"914EDECCC91886232483215450828200882112486432101A9013B3006CB81BCC",
            INIT_RAM_01 => X"42EE1F212A313100D8C12AB0CCF3C44C81F1FD3F197074BB8FF0FF0505331451",
            INIT_RAM_02 => X"10CCE9331DD67FBD34EB31DD61DD6DCDFDCDFD5CD7DD1D8D54B9D73B31931D50",
            INIT_RAM_03 => X"7F0239313215221520EB30C553C8D263CE347223C911C831DCE70CC5BC433167",
            INIT_RAM_04 => X"E60D1136016D5D5D6F010A6C373890AF015F014A466464AF012B27D272BF017D",
            INIT_RAM_05 => X"FC08C920DCE498C4C5D1C7C03DB462C4093C53480920BFBD260017471F373F48",
            INIT_RAM_06 => X"400CE60C30BC05B57575BC0899B0DCE2541C066D505D6BC050B0660610BC05F5",
            INIT_RAM_07 => X"482CD9B2082CDC8ACA20B500372064356754447AAE0BD9A1F1441CC1C58057C0",
            INIT_RAM_08 => X"A85111D999A1444746549525457245104105125D52649C2CDA2C808144477667",
            INIT_RAM_09 => X"1749104426735C51C609914152CA7842645D25755C74C9D75852449138AC8187",
            INIT_RAM_0A => X"4519A07182558DD15132576473343533834173560018101C90D9941872060705",
            INIT_RAM_0B => X"88D167088916732341160550910662878682894051428AEF306C215499A05171",
            INIT_RAM_0C => X"AD95A2C71851046589484D330AA91A084E8A9442B19B73646AAA882C669C190C",
            INIT_RAM_0D => X"25544616CA1B61B5DB794085561A755CCC49433304D182449D083A003563548C",
            INIT_RAM_0E => X"1112710A81111720A9111174572531124805D141D7314041848408CB5B4B296D",
            INIT_RAM_0F => X"C9D12106340C171CC1898909514CD281D1D810736710A81110710A81113710A8",
            INIT_RAM_10 => X"7074A0CC1A388205C0913B34D1AC9C58217258AE600381504114180E4D928184",
            INIT_RAM_11 => X"0C5536D58640966084642E994325C8008C55215405501922640990C1294281D2",
            INIT_RAM_12 => X"73544655491913665604260416240566448D1004D99CD4494485574B74654989",
            INIT_RAM_13 => X"409150404410C01F0411351251A18196D19595D1915504095509586065B05506",
            INIT_RAM_14 => X"915832130508154104081432424366055298D9A898D90D9EC1B34CD9C145411D",
            INIT_RAM_15 => X"D15989CD45C11741458455710C71861451041289C51710C718614510412853B3",
            INIT_RAM_16 => X"310050418706656474ED2914DB65205252160C7125855D173345563624274540",
            INIT_RAM_17 => X"981D09906A091850D6009901D89986A89181995DD13606902E30548080141220",
            INIT_RAM_18 => X"6287872614691514453A34634364005D582470448A0404A851373137281D6809",
            INIT_RAM_19 => X"49008840909964814B4A4D19951160CAA690672349125624237392424A01DD26",
            INIT_RAM_1A => X"621505224C38C2370A5A9942300F54E64B45646419262708884015085925D191",
            INIT_RAM_1B => X"632DA5020604196081430A141A60814154418173648A516C2442637A54CBAC9C",
            INIT_RAM_1C => X"349AC8C0664475B0B2889825947246D95D9D0D2680087DE0959E215669498996",
            INIT_RAM_1D => X"64174158C112D905D0572615043407775A4549D58A11EC912182637840505132",
            INIT_RAM_1E => X"C81C5801F401ACD49D5ACD90E0D5D150508AC10845445990590541DD9923660B",
            INIT_RAM_1F => X"7A2451D9D1CA46042360627B234989ECD2696431442012314345C0470C8137B0",
            INIT_RAM_20 => X"3606342435415D51256055354C99ED50DD895C5959E99D58D123409E4880B6A4",
            INIT_RAM_21 => X"5846140744209370253448814DEB773454435411676459C50458191911A1419D",
            INIT_RAM_22 => X"431C61851441048C8D27A205792C61441D2203185107144188C3411044054527",
            INIT_RAM_23 => X"8802120380DD05B44204CD363600420B24431C61851441048431C61851441048",
            INIT_RAM_24 => X"A851511113564536599374851511113572B2762599370C1930426160C0DD801D",
            INIT_RAM_25 => X"98805D4051515110672B276269876662673422A1A0A066463669876662643740",
            INIT_RAM_26 => X"19C96699B66191745746440365374664B75275BBB8235B383A00C98818001800",
            INIT_RAM_27 => X"2000016184581501981628A610546141445754410409051019D5CD5819090910",
            INIT_RAM_28 => X"44E820524704B5D34342A919CA7841A587754415161D0800009200002880000B",
            INIT_RAM_29 => X"540035450B3D625595288041004D00C16C8458820446243DC3020449581019D0",
            INIT_RAM_2A => X"41CD9819C5DD159181D1011589189890990151644D000489DF49F6A436010135",
            INIT_RAM_2B => X"0989250874344DC620B0030000ACC080C08CC051168005364354191913560652",
            INIT_RAM_2C => X"51B299010101922932060678663406068A4141945A39059A163641564121C950",
            INIT_RAM_2D => X"312019E512A18D86D1C5C92654756152D661819A400011524968D288A5251490",
            INIT_RAM_2E => X"0D2230F2333670D2290A89E13072461726354919100889D9185D105D01005259",
            INIT_RAM_2F => X"27365B00672066272322205607064050643499D963549C08058910509C1512C3",
            INIT_RAM_30 => X"A8C2053048C10305C531624140AA258DD50150981585D200C00D2200F2300228",
            INIT_RAM_31 => X"49649A308C902452525410C214C96352665925929D364645C51C04D927592592",
            INIT_RAM_32 => X"C1A88814966080941660805D500225666644090950022592592A450D24649902",
            INIT_RAM_33 => X"24261424225440671549445619D19100994DD191000900080C129062049A8881",
            INIT_RAM_34 => X"017D42267154DD181092420508604D8098989035012501264604260424226646",
            INIT_RAM_35 => X"0160C5CD06274458314341C5D4552009D5049832434181D2260C94D070752648",
            INIT_RAM_36 => X"00AAA00AAA000000080200AAA000000AAAA0AAAA0AAAA0AAAA0AAAA014664242",
            INIT_RAM_37 => X"830080808080AAAAA8000005800000AAFBBBB00000A220AAA00AAA00AAA00AAA",
            INIT_RAM_38 => X"5500015500095580208200000000030007BC71A3852CC0300CC0030248A0F0E3",
            INIT_RAM_39 => X"D7004A00963C6FC8D714489CE414144440282D88C11414444001550001550001",
            INIT_RAM_3A => X"0AAA0A2644C6C6C222222222222222222223332279CC4933333CD0244F3C6FC8",
            INIT_RAM_3B => X"7EC78F303302211122CB8844D84E4E943E90E43B8E43B8D03E0D03E228002800",
            INIT_RAM_3C => X"A000A241DA41E4D5C95057140C18F62E38F60C18F631464471BF0D00000000FC",
            INIT_RAM_3D => X"FF3FFF3FE83FFDCA140113535C96054818D1884A1F0DD18801C44D70D4B72A40",
            INIT_RAM_3E => X"80820048021003022A160041FFFFD10995DAB90CC330D8793D8A83E43FD8093F",
            INIT_RAM_3F => X"327010069ABABC000F5D16880108542A285502169002A0160042900290206021"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"92C7EF589918C63264C6328000C28314CC30424CA863052AA141D102FCA0B001",
            INIT_RAM_01 => X"A3BB191A370323281E0A1DD308EEC44072E199372EE284EEC660770A0C260CE1",
            INIT_RAM_02 => X"240C95001993015C644782B1F2B1FCC44CC44C8C41192E0C84100808644027B2",
            INIT_RAM_03 => X"3C03F5FC333B3333305520855044D370453483110D61C402201600C548937156",
            INIT_RAM_04 => X"25B234CC071F1F1F1C07B232C9C9CB2C070C07414554541C077074F7470C073F",
            INIT_RAM_05 => X"F00F151B272453305CF3CF0B40C49313480CB00B5511CAC114D273CF3C13C00B",
            INIT_RAM_06 => X"ED8725B21DB01C7C7C7C701B84CB272712E01C0F202F0301CB4B65B65FB01CFC",
            INIT_RAM_07 => X"761CE871861CEC89C518B8243A026024A7B4B4A61588F102E34C30C8F301C301",
            INIT_RAM_08 => X"10DADA9E92434B4A4A4BF2FC5862CD30F34C301A1FFBFC9CE51C60037B4A7A78",
            INIT_RAM_09 => X"1F87A2EB04714C000203E0C3328B70A0C83A2C8761CA4AF3C1F5C9327DF4ABDF",
            INIT_RAM_0A => X"492653B250A5B529294E4974A3383B0143B14397332864DCDC59261741278C0F",
            INIT_RAM_0B => X"89724E089B24C125D32407307A2EA20D0AFCC1633CF3B3C8015C12C8321022F2",
            INIT_RAM_0C => X"B7FF324F3CF3CC8781CC05C14AA8343709098C89737B93A26AA9361CDE8C2800",
            INIT_RAM_0D => X"0FCAFF798B3EF3CF7DE1C4BBCFB8FC90008260022772A90419801732DFAFCAA4",
            INIT_RAM_0E => X"3080402A83080402A830904855229B648A82A843EC3740C2BA0E104BBFE12DF3",
            INIT_RAM_0F => X"7912110537F05CF8098DC249F0F05D0D52542CC38402A83081402A83080402A8",
            INIT_RAM_10 => X"D14870B0573FD135C41204041218DC1A0080709DCE235724FF4FF80D42103047",
            INIT_RAM_11 => X"48151C720CA218821DA69592AC26B44AA861AD468154659E568598DB2900C2D3",
            INIT_RAM_12 => X"6274B648C5257C5849290B1909092549595B24A3E48C9FA9FAA649694A55620E",
            INIT_RAM_13 => X"4111609178F0085E00D7077877AE0ED952529992D2D244A4B30BBB83B671953A",
            INIT_RAM_14 => X"60582290090852C54058241250A196185298E9505461CE90455140211148C521",
            INIT_RAM_15 => X"12128949C9C904A0498892C124E34E34E34E3042092E124D34D34D34D3042040",
            INIT_RAM_16 => X"9111A4C1BC34B484A0482104B1C93229F0ECF4C22641212320484A2626084808",
            INIT_RAM_17 => X"AC694A54DD0DA4A8ED045A8A9CA54DD8D242D5DE16B81A11280185044A693312",
            INIT_RAM_18 => X"A20C091708552F0CC524249273845D35209490A00548805C292B101514D6D445",
            INIT_RAM_19 => X"460D80C4A86D9488A7C081212552C34D99E05C108520C8392971517085C2560F",
            INIT_RAM_1A => X"D10BBE1085D76E0A026667C312A5CA5E024BA66A968809377649C2B7330D6D29",
            INIT_RAM_1B => X"22298305D75C10929244D34C10929262649252738489F2C2E4A28242486D75FB",
            INIT_RAM_1C => X"97E0000147487A52CF0418B6780340DD99920F3F008B6F0887E0BE5FEDA606D9",
            INIT_RAM_1D => X"4A4F57200611D293D5CA18181B0834A5A644CDD68832002DD362824380D82D12",
            INIT_RAM_1E => X"4ACAE30C9EB3A8E099694E9C949D2D589041013448C86D293D5C8D2DD290B707",
            INIT_RAM_1F => X"A5249219924A48092290824021F349049CED96D047DCD30042498B0B04ACCF30",
            INIT_RAM_20 => X"981919046C9BD2DB3490B40B60D2DD642D0EDC2DDE1D2D6C1121E4900044A666",
            INIT_RAM_21 => X"C3DD15144A115047530484908701F9454CC6C9B4D49652026D30256591409B12",
            INIT_RAM_22 => X"4930D30D30D30C0487CD228CB028E38E3E028934D34C30C380C6D726E85C935E",
            INIT_RAM_23 => X"80A282802CEECE76543A42B735266712144A34E34E34E34C04934D34D34D34C0",
            INIT_RAM_24 => X"10D2DDAD83544A0855504F4D2DDADB35405049055504BCA2C1B0808709DD0991",
            INIT_RAM_25 => X"24442D84D2DD2DB0643534936775A6A2A4050343536067480B6777A6A2A704F8",
            INIT_RAM_26 => X"C8C1C8721C879B4B566A4A28A2264A66A66A66957102781515208A04A4446C84",
            INIT_RAM_27 => X"213224A56464524618595019C8948091549449C532C282C019D58D5419C10D22",
            INIT_RAM_28 => X"E4C0C4994830A7EA62B2A9294A4377B667A49C56199E0C4489B2112268C4C899",
            INIT_RAM_29 => X"18892E818B2389115EE7609B209B808D9884928A4C88150F880008A5202825E4",
            INIT_RAM_2A => X"690924290299D29A8D1229920E949C24658619DA6984A66899E99EA0892E8B2E",
            INIT_RAM_2B => X"26063A77790B4E01174DF6C0C993099F099B09291902293846C9B999B2492A42",
            INIT_RAM_2C => X"D2629242428A932A00092A4248090A194082021C650216642518421FADBE0D91",
            INIT_RAM_2D => X"142469012242495D3289C924A4A497293CEE0EDD4040109361989348934D2CD4",
            INIT_RAM_2E => X"7710175101085741298AA900015049042826816DEB1C4DE96819682986CC1947",
            INIT_RAM_2F => X"143A42029400950B302021861A395293941F39E98E48994089422C2498613261",
            INIT_RAM_30 => X"B60709C0AB02AC2AF9C2609080A92639924A182C218290126237102351023916",
            INIT_RAM_31 => X"A9CA5981C45CA4805168A30727058E51587AB7AA5E6E4A6AB9240CE8B672A72A",
            INIT_RAM_32 => X"C650986CA1149C2C21149C29A247057664A381C5A24707AB7AAA4A39FACA59CF",
            INIT_RAM_33 => X"0A260A2600448B23376B5B44359A928A2889A292AF02448849B29A8240E5098A",
            INIT_RAM_34 => X"91628125514499A064A092024A425B495458146D26152605481A262A26035448",
            INIT_RAM_35 => X"0142018EEA0A48108153BA0298511249BA04508243BA8693242058EE82A62544",
            INIT_RAM_36 => X"4BFFFEBFFFEB802EBE0BEBFFFE00A80E757EFEAFEFFFFED5FFEFFD5E24A4A050",
            INIT_RAM_37 => X"FBFBF7B37F3BF144195555D01E3D559122EA6C2B2C10201FFE15FFEBFF40BFF5",
            INIT_RAM_38 => X"EA800C258006AA4004440000000003040FBE9980B0E0FDFFEFFD7B5C844CFFFB",
            INIT_RAM_39 => X"4300370C433C37CC4300F8A45714A3482B14A3482B14A3482B0960C00965800A",
            INIT_RAM_3A => X"FA500FE98C2231867EF4444474555444445CECD05B00FAFCDE14CCF44F3C37CC",
            INIT_RAM_3B => X"3FE2FFC23C0801403E0EA050FA5003E97E90FF3E8FA3D4D4300C03F2FC16ABFF",
            INIT_RAM_3C => X"AA50FE9D2591721C418C71230D14040D04040D04040A081089302683A453AB5C",
            INIT_RAM_3D => X"FF3FFF3FFF3D40CF282276909CCF46F44E9244DB2F270244829D8D81A847330F",
            INIT_RAM_3E => X"29085921148A575480806A1455AA9FF6AD7D7BC38F1C386ADFF7BEAA9DBC903F",
            INIT_RAM_3F => X"E814800C0000000005500012A892014002005840066804805628049409480580"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"01068A44400040110041114000400100442000044411001010019102E773C021",
            INIT_RAM_01 => X"22AA29282A0222281A082A9208AA8880A0A29A2608A208AA8660660504110410",
            INIT_RAM_02 => X"0408AA002AA88006A816015011501641064106A4142A0806A805502A655C0622",
            INIT_RAM_03 => X"010905053104111110692F8960B8A2A0BA28022E0A428BC00026308988126266",
            INIT_RAM_04 => X"0001120504000000010500040004C01104210611111111210501011010110400",
            INIT_RAM_05 => X"04242440000148141000044020010048000000002440000052004000110908C4",
            INIT_RAM_06 => X"4054110150441000000004141010001320141000000000410050110110441000",
            INIT_RAM_07 => X"038E2B38238EE7D0E38EB9DBF24D2CA0A2A0A080A2D0D122DB6DBACA49410841",
            INIT_RAM_08 => X"828A8286820A2A0A0A19004800A48614E185320E2439298E238E088A0A0A1A08",
            INIT_RAM_09 => X"5194651BE2A49649A798261849D0589539465084210BD218E9043942410D296D",
            INIT_RAM_0A => X"0A488C248C0840200200080084D2F1489E3C2F09D26D21232120218438C8E394",
            INIT_RAM_0B => X"D01620AD09622B40492294494253B4148AC40835049010E18682C5094EAF259C",
            INIT_RAM_0C => X"095CA4141041048008ED0104A00BA86A6A1AB7D4393B9F2D0000038E4EB12B2B",
            INIT_RAM_0D => X"600901F29096C14C97C8ED051572018E10161840484422FD82108A4A0481492D",
            INIT_RAM_0E => X"1308B40031308B40031308180B42CD22501164D44C5115912B1C8AD014CB425B",
            INIT_RAM_0F => X"4002695848436202323270322903603240616494AB40031308B40031308B4003",
            INIT_RAM_10 => X"859A7903A68C08E9674290DA42692963942D8A22106990A41741772692AA8880",
            INIT_RAM_11 => X"1312640214B41489108BA81220CCC12A1103308F312703208F312BE6C322F6C5",
            INIT_RAM_12 => X"9DA2A209280A61090848404841486A0A0A902D2579B285C85E2A0A921A20923E",
            INIT_RAM_13 => X"68868C8E8209ADA1A3A6907907821076C6C244424242D0205729F8841D840970",
            INIT_RAM_14 => X"AD9AA44841A1D23D10F50694C50E0C70FC3FE313312A3E325A59E12A4A09E828",
            INIT_RAM_15 => X"4E4216F656F2908D09A1422A6143143143143290F420A614314314314329090D",
            INIT_RAM_16 => X"8D4CD0C9828280908E23A959800B4A24D2A10638DDA424E595390859D949392D",
            INIT_RAM_17 => X"2103583FCEBCEBC96CD21AD03D03FCC3C290C3CEC67840CB42870CAD02343A40",
            INIT_RAM_18 => X"B41489594264209216A8E08E84AA410C23B0851A1E125AE52CC0CABBFAC2E121",
            INIT_RAM_19 => X"B024212301076D28934AA42424421867760A638424660848458D359424564260",
            INIT_RAM_1A => X"084080842000004189D9582A40A14916CA09A18B42D8526222F6926A5F2828A4",
            INIT_RAM_1B => X"7B4D25A00003B98E87A20823B98E879DB08787B4AAD0D22520B458CA0A000008",
            INIT_RAM_1C => X"05F2210A664A49B420E1A19D8668A24424429658E2D35F6D34B293C2E4E21076",
            INIT_RAM_1D => X"094290AB10EE82D0A429C0C2C0C160A0AA31288AD052290AAA3458C827A50AB4",
            INIT_RAM_1E => X"D094C8A96C832707A82AF0A183A86827AB261EAB0921C8250A42A82882ED2A72",
            INIT_RAM_1F => X"B87A8A8CC29068C84F8C14CB465F132DC3E7652790C3E5879FA8D248AD095C8A",
            INIT_RAM_20 => X"D860587A4290426650861949B54244210650650642A42421AB46513221213B31",
            INIT_RAM_21 => X"D06C79F3084BAF90A7A0AD0F1B200A221214290420AB825A410B482ADE2690C2",
            INIT_RAM_22 => X"9850C50C50C50CAD197CB4448B4451451228991451451C710AE410250A4290E6",
            INIT_RAM_23 => X"30B4044887024982A0C93280C1DA958BEA9811C11C11C11CA9811C11C11C11CA",
            INIT_RAM_24 => X"A1C2ECAE5F0A094288A6942C2ECAECF09616086802694707043C1C1C16203680",
            INIT_RAM_25 => X"05210292C2EC2ECC0971708783B080860B6A4B87878C0B09438B3182840A6942",
            INIT_RAM_26 => X"9B2108421084261A0A1A0B446CA28A2921F21FAA3849B36869D2522101210121",
            INIT_RAM_27 => X"F078D88892DA4210B3B6B1B6D8B08487B0A309A4B5D030F202C2BC21025A9EB4",
            INIT_RAM_28 => X"D2A1236D09490438CF8C010370CB139DA3B09A4296601C1A360F068D87C1E362",
            INIT_RAM_29 => X"A2D1D52AD0D52438311DFD02850A12176D1489100518D84F3441512423607620",
            INIT_RAM_2A => X"965421065064424A1682A64212633103C358340DA3B211BB86E86E054952D0D5",
            INIT_RAM_2B => X"A2101DAE7842EE3D8C10800A1604360836003624B62AC0CAA4190466E508E195",
            INIT_RAM_2C => X"6A24121834303A4684D0C0C908487049A218FCB52688EDA0E84AA2D2EB5314C4",
            INIT_RAM_2D => X"E843032C29052400021616909090802407E2107B98348C0EEB6D692D01242167",
            INIT_RAM_2E => X"07849048494A905843901327868F087B458DA1ADE45651E121312103585C38FB",
            INIT_RAM_2F => X"CE78CBD40CE70C484C8C870D4BF0E48F0E65F123504A11212810212135838449",
            INIT_RAM_30 => X"0D15A50618144041C506842C25004D43121C3121C310394A4987849848498684",
            INIT_RAM_31 => X"EF6EFF456B3145B5F5DA543594135044585F35F8D25B4849C861290B8E1F21F8",
            INIT_RAM_32 => X"1611A1052331A10B2111A103691584B48498575769958573578069412E6EFD12",
            INIT_RAM_33 => X"4BCC48CC5C4ED26CA2921A0C538686D15B286286542E161A3A4C3A84E1631A10",
            INIT_RAM_34 => X"0C1728C0CC0E312121048452118596D679797358D8DDD9DD484BCC48CCDF4D48",
            INIT_RAM_35 => X"9434313C6D40E71D0C2F1BD03503B4305CA31D0C1F135039C3431BC4F40DC0ED",
            INIT_RAM_36 => X"0FD07FFF0FFFFAFFFFAFFFFFFF00A80E757FFEAFFFEAFFD5FFFFFD5FA2848E84",
            INIT_RAM_37 => X"77C84400C8843E4E4CE4E4800CFEFEE095D9517F7C00000AFF00AFFFFA00FFA0",
            INIT_RAM_38 => X"C9000C90C002AA001405000000000303900000000500E33D7FF48F200000FBD7",
            INIT_RAM_39 => X"2828908428149044282854545414184480141844801418448006B9000C30C000",
            INIT_RAM_3A => X"00000FF34A43E9033BB10F903D5E5D6A8E921101558A55447600745CE4149044",
            INIT_RAM_3B => X"1073CFFE803A81543FFAAA5500000955400255956559565495254903FC000000",
            INIT_RAM_3C => X"0000FFFBAAA2AAAA8EEBAA3ACB18FBFA18FBCB18FBD54BB822EB2A9400540307",
            INIT_RAM_3D => X"FF00003FF70000CA0012EEA038BBCCF8FBF0F0BC353F00F042BB8B03A4B92EC0",
            INIT_RAM_3E => X"841A510848016A88C8D0C1617FFFC1159A9D1B8CC3309C1B49F0AA94EBFD003F",
            INIT_RAM_3F => X"14102CE16AABFDFA50000000604004802900220215400410A800044005A52104"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C020001114451144511447FFF70FCC7D12CC45131144C347C4C5D9BE34603FAA",
            INIT_RAM_01 => X"C44043884CB8405D401D4106010114941614104C410481101140443F700C0300",
            INIT_RAM_02 => X"00100C0C00000C002002046464646313131310500C0C4C410000000100204044",
            INIT_RAM_03 => X"20002020344C4C4C440C0300C090040050000009000000C0C180210200040050",
            INIT_RAM_04 => X"8CC80D20002320232000C8732023308C002000C8C8CC8C8C00C8C8CC8C8C0020",
            INIT_RAM_05 => X"8000930C808C34808032030891CC873488208208930020230D2200C80C2024F0",
            INIT_RAM_06 => X"32008CC80230008C808C8003DDCC808CDFC00020202020000F0C8CC8C0300080",
            INIT_RAM_07 => X"D820028248200CCE08209040FC00888A8B89888BA3FCE2E2D30D38C808000800",
            INIT_RAM_08 => X"A022222A2A808888A88B20C880BF082C820B222C2CB32FE0082090889888A88A",
            INIT_RAM_09 => X"C8B2EC8BEE8CA8A248322CB282CC889C8B22C882A0A9FCE3AB2CBB2ACB2CCAB8",
            INIT_RAM_0A => X"8BCCCCFCC8CA122212B48888BCFCEC8C8FFFFFF8F023232323222B21B0CA0B32",
            INIT_RAM_0B => X"CC6A2B1CC2A2B33182A272832EC8B3388B5C8BBF3CB2F2EA0EA43CAB22B30CBC",
            INIT_RAM_0C => X"C688BF1820820A8E8A83384C95524CCC93332CC382E80FC895561820BA23C22C",
            INIT_RAM_0D => X"23843A62CCE88698288A8CCE1A621AAC333AB0CCC8E8B2FFB2334FCF286184BC",
            INIT_RAM_0E => X"6E81BCEFC2E81BCEFC2E839B9B330EE2CEB211B280E02CB20C3889CC298B31A6",
            INIT_RAM_0F => X"D22234C9CA532B6C32323332A213633269630C8C2BCEFCEE81BCEFCAE81BCEFC",
            INIT_RAM_10 => X"9CAC9293AB21A0EA8F224CC9263B2B290CCCA8B397CDF22CAECAA376F0A48BFA",
            INIT_RAM_11 => X"2376C8E23872384838D8BAA6942A5F3E2237A5D8276237A5D82763880A2230AC",
            INIT_RAM_12 => X"9DA9A98A0686958988C8CCC8CCC8EA8AAAF22C8A622228B28A2884489889420E",
            INIT_RAM_13 => X"B08D8C8DA482CFAA13A919AD9A822322A2A266626662F3F1AA2AA888C89ED9DD",
            INIT_RAM_14 => X"9CA86390CEC3223233233B0289CAD8DD80A30AB3A30A74A27682C30AA18A8626",
            INIT_RAM_15 => X"222232323232489C8A8322B3F192192192192233322B3F1921921921922334CC",
            INIT_RAM_16 => X"C88C308A9B0B8888A4690BCB238BCF1022296CB0C892222A0C8888C8CBC88A83",
            INIT_RAM_17 => X"E336336E9B3B2233E333623362F6E8B7BE2FA6AE2538CE273A0DD89F3F0827CF",
            INIT_RAM_18 => X"B33888C8CD326A20325CD88D8C29CB2A13A88CC23B3332B330CC8CA8E9223336",
            INIT_RAM_19 => X"2326232232322F3C40889262222292C332913B0CD22C88C890BCFC8CD3F222C8",
            INIT_RAM_1A => X"A0CE5A0CD38E38CC8888CA87CFF38438888E88E823088FCCCF33210CA62222E2",
            INIT_RAM_1B => X"83F2A810820AAA8E8E90820AAA8E8E8CA88ECE8C29CC222858B391898938E3A5",
            INIT_RAM_1C => X"EA222234888888BF9640A388A4924222222272CA42CCAA2CD9A2A266A8A22322",
            INIT_RAM_1D => X"84CAB22373ABA332AC89CDCCCCCCE8A8AEAA0AA2CCE2233AB6F3918A43A33A73",
            INIT_RAM_1E => X"CE2A8892AA92E333AA2B33A0B3A26267A6D33A6EAA033A132AC89A2AA30CE8EE",
            INIT_RAM_1F => X"ACE96AAAA2CE88C8CE0EC28B3CA20A23B5A2297EA1B3A80E8E9AC8889CE29889",
            INIT_RAM_20 => X"28DCE8E9C8B2A1A3E88CE8CE83A2BA233A33A33AA2BA2A23A73CA0A223226AE8",
            INIT_RAM_21 => X"A188E8EA88CE8EA97A189CCFF2238A9AA07C8B2CA8E8A232CB233A3A0EFCB2A3",
            INIT_RAM_22 => X"FC6486486486489CF288B3C89BFCB2CB2226FD249249208289ECB22CA9C8B2B8",
            INIT_RAM_23 => X"3373C9089310C89998C23090DCC18B0B19FD2192192192189FD2192192192189",
            INIT_RAM_24 => X"732122120CD988CD9DCDA122322320CD8DCD88D9DCDA173A4CCCCCED30663062",
            INIT_RAM_25 => X"332336322322320DD8CCC88C9CC89B8CD8D9C8CCCCCDD888CC9CCB988FD8DA12",
            INIT_RAM_26 => X"222384E1384E609898988B24888848848AACAA9DB8CEAFDCD8E2322333233323",
            INIT_RAM_27 => X"CCCCC099888922332322333228A88C8EA89A8A464A3333226626F36376767272",
            INIT_RAM_28 => X"8223632D8ADCD9E98C095A8A028AA688ABA8A4622201FBFBF00CCECC03B33300",
            INIT_RAM_29 => X"62C8EF26CCEF2266694CFEC64EC233322CD88BCB0A08D8CE38CCCC1623045500",
            INIT_RAM_2A => X"463A227A33AAA2A23AA242223020A3B376376270A63308822BB2BA220882C8EF",
            INIT_RAM_2B => X"E223089DB8CD9E374E38E389300E300E300E30222224CCC29C8B2A7A3E888E8E",
            INIT_RAM_2C => X"65B3A2333333A7390CCCCE8988C8ACCA422FEF232908C89CD8C29266A522088C",
            INIT_RAM_2D => X"ED077A2A25CDD618623636589B98861069A22323FB374CCCA22365DCC6262363",
            INIT_RAM_2E => X"9A0CE9B0CCC2A9B00A254A290E8E88EA391ACA6660AC3AEA63662336373769AC",
            INIT_RAM_2F => X"E8D28AFEDBFDDBCBCCCCCDDBCADDBCBDD9CA2A0A9589A62326008323A37673A2",
            INIT_RAM_30 => X"AC2B184CED33B4CE184D8CCCD2542A5662376323763367CFA21A0CE1B0CE182C",
            INIT_RAM_31 => X"A59A670AC3A228BEBEAC252B213A958EAAA2DA2860C98A8A16633332A8A2CA28",
            INIT_RAM_32 => X"327363332773633327736336B02B2999A8A93A3AB02B2A6DA68A8A566A9A6636",
            INIT_RAM_33 => X"CB28C8288ED9C88888489898E62622C9222292211222363A3680A88293273633",
            INIT_RAM_34 => X"8DEE25DD8DD96623224C8932248C32F0A3A3A0C8C0E8C0EA88CB28C8288DDA88",
            INIT_RAM_35 => X"C9FF273F8BCD927FC9CFE2F362767237B8967FC9DFE2F3659FF277F8BCD89D9C",
            INIT_RAM_36 => X"4100041C0341FFF41FFF41FFF400000EFFF4FFFF4FEAF4FFFF4FFFF45AA8828C",
            INIT_RAM_37 => X"9755555511112AA553AA550006565560EA66640104B200BFF41FFF41FFE01FFF",
            INIT_RAM_38 => X"50000501000C00C024C600040C0C6F00600000000000E97A4CEA53900000F8E7",
            INIT_RAM_39 => X"9614E948BD004A0096000000000000000000000000000000000AAA8001450000",
            INIT_RAM_3A => X"5555500EA554000CE0256A96E966A59565A66660000000AA9928C88892004A00",
            INIT_RAM_3B => X"B83FC3FFFFEAA955400000000000000000015555555555545515455001555555",
            INIT_RAM_3C => X"555500AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8000000229",
            INIT_RAM_3D => X"FF28003FFF2AAACB2DD0000018500500C436011443400A012C00150451108215",
            INIT_RAM_3E => X"018000A112880012E2C5E804266ABFED5AFAF7870E3C70D5BFEF7AAA5FFC003F",
            INIT_RAM_3F => X"65500870000001000000555A0A12612680994860402992850229521680008091"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_3_AD_i
        );

end Behavioral; --Gowin_pROM_cart
