--
--Written by GowinSynthesis
--Tool Version "V1.9.9.03 (64-bit)"
--Mon Jul  8 15:35:15 2024

--Source file index table:
--file0 "\C:/Users/stefa/Documents/tang_nano_20k_c64/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/Users/stefa/Documents/tang_nano_20k_c64/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.9.03_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.9.03_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
EqpCJ1Ww4Pd49B2vVASAo8LpiKKOyOr3fTQtoLEopzYBtsWzW9bwJBFufjYHFtUn8GTtPZPMO28v
8B5rUJs4Hd9uLl1OBi0kSgzbjz0PQjZvvBaG3FrvJm5WkEEgTZf6h/XYErPHf6a9ePw1mQcK/w0V
Tmn92XFVjoSysDTE2lJd41btgDYM6X3vHBOaUt+NLuypAHF27Vg6/a/ukPi+VDsF926BOYJWViP6
U+svy8MhF74v+ClimO5vWuc31+6F3fQYnS+kNuW+etjyU2ZvlGD7zxUmuTqySt4hpy7pKWiCeO8I
zxJ03vHaeP2blj3EFD5TOylCkKAc+X9MKyoI2g==

`protect encoding=(enctype="base64", line_length=76, bytes=12560)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
KE6eVmjzw+3Qdz2naZJ5i89PLu3/QvnIlM7WqGHGwcxE/On9Akyt/94easmIa3RDkNz1H8r9GmR+
j0KfuHfEo5pgFd/SGAAnW5H3d2pS7SOMIBblzCQOVHx23/UaTwEbEcaDlcPjhv2W1ypk9efApsTf
ktI4B+DhlVWpOMqNXPFF01PEPccXvjpDBsfrfy/gpTTluei6uVK+VGENv0br1mey9wTajKvP6hAE
gJzb0NcqBeLR5OBzTm+cYnDpax4Rz7VnfEhiso14/vBxsZ7xUv7ce6jM5oqeqlyCjmOSmRKa/OSR
wTqzf8ejDfpUCzlTbGlAOmOtio8qCzcDx5O//mPTJr6Ud0iJF2ae1s6p2hJIKNNyb92S2zP3dK98
mSXLO4wFUH+DOuikNPGdOF72YZ5fv3CnN3LuTHKxb1yEH6Kqhcd6JOKFPudnyDPctKFV1dSMJbAT
/wTbcwTaUm6vwMQTYL3StlFK9rwiMoli+aLyoJdrivdMl+3lvhlLGZpuGxCz4Hs6KN9a9kY+yyyI
oqgxVBHjUqL40ONSox6w30mg3xV8GcYaXljNdSRp2bo8Xyi2mn9YWC31buSdBsTUoJAOvkxvg1gw
MVCUXakREqhzxC1TbKXbhdkt1pXkomuS0K5lHEElRUiU4iIGqdbtdcUqeW+RosjJf/9P3DaOF5iE
zmeO0czx8gu0qOhLObzvRyXjN7o3sbz3Z1qqSCzRULa37XZhuuZLtKPASK9e3707gpDi6GAARp3H
SMuS/rjOuaG/i3rDUlhACvAXL2wArT8GOm1g+XM0npFvzcG5CjW/M6ti85yazylNk9GhEV3QKVM7
C3T/4MJ7ZjR1li50yl3kZRooDME8Oj0K91oMOhEm2BxRckK0/CaKDIQlEBVHxcM0Wa4Oa0xLt8jt
JEzf5xcyWKVzceIyvBQ+VuOSqWDYclNHYFBf/ZOCUQcaFfcXDxjaHgT2Ris7mDuw7iHWd4IM06z8
5t/xvljW++/xvOufXuNcxcY6DFY8D9hSsdL7/H5FIZK9TKCXKYgU1RsNbhTq/mQE7U/M2Nn972a2
F4iXB286dHucbzBwjHRzAVJi6QsbAQRzP5yAJ2dKTsJTGvl5NBxHCtotyBsj8S+5eg/RdDvgzy5B
HNSpyQCbNIR+oi/UFDIZicMzhIcHQwOrjG3l6+vnU3n9nJUmRY7E1JVU07xDL+qhhd2v8S0F9/oI
8fNGxf76orP7rQxcBCAWk9HCewWDxqtE4D1YvZO4HKyVMgdvW4pVkzs+BpH4qGpuizZS800qrmpa
mrJpk/yBU8qUO0dNE2dB6+R4hA/YI+unPhgisaQCf3iSVt9ICRsTedj0ApJ1yND7XwdgclaUS5Nv
fCoI3A2boHfsMSrKfT4gUpiQnnOvd7HD1L32Nu/xJz/SayL72SA8kLPkZZRJHOT3WRSWI2bPiU7h
2mrGKDC6c06N0Q4RzatI5JRcNYCui51pQNRS1QOW5y7VjrppIYzRYZx/rhPxJhh9IOL2eIF6cSoG
z7Bt7YwJOvopgZIlh/SCD9Mpxd9v8dcX47zhH5OwQo5JVrIOFHg3peUHyPFdjmmwM/5ls8z/AwoV
0GwJ8GoDEdM5RS+yXciBC5Qbq1dJz6urCqLZgJ/b5hceEjygW+a6ZoNFXqNIyLy/4jrm7f/XL9hM
ff5gLKX3bPxW5GVQkNM4IkSb/ut2hAzazLRrYmPjym1sgQeKR8t22wAnMClnhxY9EpdT2hwR2EBT
jcsNtiwImTp2qRHMjpgdygPiJQyI9dOcVAJk2F4Yq89aaq+ugux2BU017/8RWJLadAbji8guIuXZ
BmLkJP5kzFdCoAYoVoEAbfPtvemu0VHv2U5Ec4/BtdaNiiAKjznNB3M5hHhRjo2Gp1fWQ+hT9cqQ
z4N+iggLkoujIjXYVIgT9RJZtIxR1UBFC4CQQ5EVzcKSUQchI5KGWdic7hGVMgXKT6lVZGpAnqtS
RUYATj45JjBMWjkE3N8X+pv2cYcuwKHGwwaGdzQErN+gmNPq5GZG68vnjOMnJA8N4GWV+yKDGi9t
M+arA+kw7JYsIiYx2VMMye0sG1bG4weIDFO8ZNXMX/IHFAy1x+RH5LxinlICPv2HCjqDFrzt9RTA
GBCfPQEJ3K38IKZpWcGCqZywbcBQLRyd+/VMWg/YzudVehDL67GXP/UAuJuddS8qqw76J2JrbU2k
ybXzFeDEVd2MAp70CmvbvtcNTHbspEDJx3bhjpIUPusMofPZZYFDclwiVZemn7L0QqVxLH6gfsRe
HT0ITrJCGWFbzL25cl1v5AfA6zANadkFi+j6N+qrBnOu+uQwWmPnftqNJ06PIpdmvW/dfrVzAFo5
qkJcpSQoeY2OX8yOf7PBi/8z9cDJVITa2S16PhgVRKYEH8qAOwcKoGTccy5BXzNyoj5M+bt+uLzx
0oWyZxgeY047IRYIX1uT+K8eemK2GXK5/Cp2xMwVSzN7YjQt0DKICuO9ZDXeZufwSoz6mrbSZz/v
My+YV4QqPMWSfsdHVO0YgivlHrir20GIj61hbe7CLzT1rqHqz7sXZ7N7UI8fB7JQtm2mBKQbU4KR
7sw/6WqF62Vj7ytDvndbp0O8U9HQhp606i8xpbejlJyoGdmS1TGqqV1rMRmmXSN9jktJznd06fHL
e1BIYGw/pwjP6IW1CVU+qWSJWoe8K/AdLTJ1NOVp8rdhpZZYdI7cNTMgP2gMAdibVFjvYCLpTRBR
VZl+niDuVutwZXE94c9iVVJ/O5a6gqT/deKSuB0gm+4FcrMi2pc9bMmK87YNI6V3ZndHdbhs1/Zv
IYi0zUZqaYXYFT6QnfFRllMGs3RQ5HsX1dI0tMgoxJOAX31BuMKFUBVbmAE87MJD3gtvXb49jn4G
Es8ZiFexdGA9UPxEXPUi7a6aehlK0QKxpDReanStP4qT01NGCcJ1jQuhlj0QRLFgIMEuajL9Tvrk
Xls3pzJoa2RdQdi8lLJn7hoE0MKarqR5heGjUM27MZB+AfOw7V2QDtMXNviWQYx91uR4+8hK0cFk
fdW7nfL71ZRUwqHBkkaiACKVtGvX2B/NQ3UrTIbLcAXBjppbSk/+Gu8R9Yp0tmkJTxkqdX9fm5FY
odOX40AcZlZqshI6UGRfMMFqxe9Qq68n9hJnPRENcaes/e71RxcF1Hu9cGDYwMOsb4JZQjAcTfxU
uJDcYH4dwwgTQE8QIzytXaYvZCEcW+XXID1w0Kdcg9y8XLUz9JdetqOkx0PnByQFbeOOing0KcF7
iB5MpNiCVqyM7UjytkS4HqRgOIGaPhg4n+tMP9kkrn5GABNbyEmCKLe66y+7OfzYZAx7ZwcRaPwI
G/+c/SwSYi3feTBv/d2Cx3De8n3esD4LsTEQ8jNK4u65K5YlYW9alNWPxDDTtw6tpKMk3ZDKBA9O
2ZURC8JcjS+/7sMEEA6OiTLKPSzWVKXFSYfDMyRvzuGekvMuU7pVykdRIMZ9vfQzSm9EZWL7O36r
cFrYT+X01pS82IT7Fsl1sHs6ZPVk92AFORw5yL+9zJTnH3ByrSFvMSaN2YOrOW8erKzWifbzdKXR
9/8sEYpO58Im9QLm3kx4HglwLrmBOH7nQs2T6GB9MO3l92jR1aV2aN0nY7Umlx6R/4slgyZIe4nr
knnSlnzM/nAIc4O/1KjMoNFp8j7X96ZnF8Mg/+uyc+YmTtag/qA9ClADfChYJDyzPrG8Hs+YsqaX
kXHQktN+ewWbjGFt95i+zO+4ul8zCD0/G6CwIi9Q0xeRLs1OwT8FjoMwo/0Rk0wnA064HuGAHO0V
JbhkUbHHwnbO5ybWU2hGhjAu79INTfhL6IQYnlYwXKGEqlZ/qU0HUPB1s7FtPA0ILXQ+vePuwh2g
u3qkbgKT8ZpWHhlFe+eqHDqS5hIEC9suw660E2QSMJ9pmloHgylPGXMO2XnwkZNVX6hGymMfA9Fe
IbIQD6/1IQradaQ6jmswNaVWeycpnZyYiZmqxqHqQYALcUvl6krsUmEOz8eMxGMrkDrYNqtmUT+a
kGf/UuF/N2xHpYXvoPjInLC7QD6bv1ul/cvADjf8FVbyryEsi4WphAPdvLF8vlLrtsWkuUWNUH7b
6TVL9kGIsIcGvXRj/txTBiOQ3W+CQRRUY5MRCPiB2qPvc63VRJV+p0Ok5xIL5Shi9zZSLpRf2Z3q
Ggsw8JGqFln2EwRieehiIwNOn/5rXLJcKJ/YdqqjiGqPeS/AtYq9PWnZlglXKiRrlyiVnZeEYPfk
mmaTgieZjligH4sJF/Z3Dn9oWW1JrwkCRQWlV+NpnnsvL4ZgnBQ29dt4Fo/pWsUHUXMCCNokA9ju
C5Qok0YRWKtRA+OQeVSwHKMhH4hSL0t09sBiICZYZU/P5VoB1qWjC6DYAQVOwf3VaF8xBpQuGEJQ
FPf7NZZMiD0S7SYgDG55RpmD+rBzGYDCX+5irbAdP6C4uBuq0AkHW/OGZOC1Um+GYQ5Ho8zqGVsD
WDOX3bACoZlRj/gdU96dBsFDRBpFvXVrxTQqW0kAHBrA4qr6OaNFQPeWymabOcEXZveH7Qv6JZFS
b07WXZ6SqsPLQnOVKkA9Qs3ib0WMm5linIZJbdFDMQD5x8nRDEY6O1ygrnZcZs+nzumU24cXuCoq
JzMm/Xp71xtydxdZNblbGAndTPhf4avT9w0vkdZaZIVGjQfCtNHnOAiV5snLfHPQNZ/R06v1AH5f
kczpXHf+dEAI8LPCy1K8JweT8mWZji3v1+p0NYjiw3ViTO5DagI2R9embg3TY0QOJgN8D0cyOIvY
+LLcxwbJaAAYXig6JqhFTqYE0zXKYJy0dgu5EnG36tFfQvXMekBHFXYSQgwepoqzmhNFYo/j+n1J
7eU8VqQX9KGWgGHjynX6c2SvjtWZCcW45mCznjrKwbp7+LWDWGPhpP94Z3B28cx11s6Hh3Xe9vpi
ofn3jwhRfqkkS5Px2N53mwxzrtXrRtgtoTNjEk/GrvId6JgufJkC+G8+307WM39Ks9it0/HbVz5e
kVRE/lQtCmENwYi1YnTsuY9Fa481eH2sFpvLACPs+neu8d8PlA/jKp79IPBqUiMJVkDDDgyv5FAU
IPkYCPNApfdrjo/kgyy9SLq23nWJ6J/3kZFVRO44Fm/ioSQa8bduV9kX/HXAuDP/5Op6XHMndAKb
aXvc/ttF/nkyaO8WPpbRsTV93iferTtS41I0fAGFv7eA6sTfIk6VQSf6JRCeUi0uJT1nulbCeJJG
+pvQf3oYGbPoRj+RD6etNfwsZE2+ws5OqVUSPmlQBpZ000KydcdNKNE5rei6fQYYS+zfbejcI/oC
PeeGmAqk1S72efxnZCrnGxUMK93dYHVirEHGM8nwcsenXJ5/wgp0S/hh1y61EPGATvjuZQ7539pB
zQFDz99aIuzLWZqUoNHcPjadGXKKh/u0DxImCF+q5w+eoG//s1siPes2eqUXI/XuJBX/i+Pd6Xs1
ISc+2rpK9h+58btkyTj6mzJvAo7LLLP2VK2mt6gbsqOMzt7omiKqBIZrJVREfNnArgnpXvUs3Nmy
ee4nz00vU2ECdkvpWTKtnrRwqdf5cVVACWkkFCU1X78O2UXwmZ4IXbpejQRwxak3iAMsGG65cPqv
PNT0//ZPgTebgDkxT2wBXEfK9tG/4FkFb6Ofxb3Qb/+pwv7QNJ5oan6pzARfvVLq4RHCkQ7+Drwf
NaK9sOkhSCQ+PtxBqRsfyLu+beiaUbUiDxQkCzRI9uTsTTs8YI5ljGeDLTwTRB9e+cixTnKP340t
mhFftvAa4a0oSYrHF5vIxpRoYn0XI14/FrLKTzKFu2fRvHdkJIGA1SNGp+o7SWDEllitrMowf+Uh
TSzTZbflLwbhTdquTcdtZq7oLf6E4UQ77DGHihMriWZ56kevdIZ/bu/BU8/OnP4lhAsLM3foOBSV
QLX71/6iUPlKOGT8CA3rO6IttsywC4LyKjRzB4Ezhyfq9JyDajYWgqTbr8zzBVjW4IWLGPR/DecJ
yQbfsX5JldMD2hqzFznlpFD7t64pf4Z2PnzuWbYGhr/0XWHWsds6acaW1OCQEKnlk4uf7Qzxd+P/
aghaqBGNOYnFyQYwgV8GwyyerwNXEIe0hm2/9wJuc1KJBqLrzzHC6g9VrKpDDg+vP7TCZU8VfIxa
RUthVZGXfHP1fHd9a8rYvydQL40InDrOkSyMQRrCcIUjSNCbAm2HTE+TQybWD+QLyQrpYrx+a4Ec
pGpNU9FCWDvM54MJb3roukwhWbNvJmpTWzatKlaYq0HNUHrUStHh8w1wyivXQe4GlbJGkyZ2cWu+
t2ebmuGikhr3CFMv+r4lV4biyrc0iIbvboJXGJbcRui9CsH86RU6DtgjRAsaNl7oYP0b3MOITnWm
bfgPksiq40THnCZMgz6ELYfkrHGiGzhSpHp1RXC50aN2AaLgRSgIC+Aml/3CVa1hV3XFn8enwaiv
ciljcyr901QRTHTEIQvRDf8YFJUKIOx+p1XkDqr4VyKEhncz8KRXE26Y7NwfAG6FbFgOXl+4YNFE
G0ezghPmcekLaGcssfeCzOA2Bca9d7pDrOljwPa/v0jIUw9fBA6o1X+zdAr16eb+WZFm84waraMH
0pAdibxySVf6UwRrFQKKfqI02AOtMs6fjI5bZRDtR6wQLxwNEhdLqR1T/7rBQqyRoKGZGwQrComP
9+G0mujU0KjswxKf9HWHtrxDQlYVmLDm9zFIRMXfRdYFw05vtS1ekAf8LaV28OfGmGeqAHIaT493
Q224v5tVaX6aeqWNTbg6Cm9EwsNihSha5W1+TffNZK3BUM/+Sx3P2gyVKW8xekF2pjmrbEL6srkc
7lvT3voW3/FqX6ODNab5IU+/U6JcnAWcSAXISSR2vpDAo/Z/Osp+fJ0M0J6IjrmqMJ+cfOv4iIAw
gn3G8x0fa+2TwOa9KeqQIZQoWFJOVlRXT+2hDZ4ndzL8lE2tLKu+lenhKbbrnD7DdXJPta/4u3HZ
+VGkqPPx2ChUz1067RFdwPOdW04miANKqkHnAqQ4mVWA7/SNJ4y5OokA+ZUvzSGP+DGzSTIMYkU9
4HHHIv2tYm08LBbEh/4b98lZceuAd/7HeoK5DbpA3WwXfAbHAlt2cePqENP9Kae7hAFkPua2bIOQ
0w1UyhLP8Sbh9kMyNwilGxNZBNi/FpTf481REkTd680XlzZFleFK6GnUH2OJXw8ryjqm0x6O4UzR
zRi7WQ2zraXBF1+davh2aVH2PVnJ5IdSECFJbkrmBxAKiHAi51LjBXIrsgpFD47SQ6P+0aIYWDjS
YLW1HSa4Ng0NOVat6firBNTyl5CQoHFv0ASIy6y34k6Ir+tY1xtuzOqthE5H5Kdd2fYLupof7dq1
ff/rDL1gnDNAIyy8Vy1HmbTaZQ9mSgOKeHmgUJus9FA1Q+TqhWkvTPTQuX6orbYLA4AvSDNki8Kg
gCAIQvrom8myffH6pw5kkL1ELnrW6wrrEgMV6srUzcYBbUEPSOgg2+pmbyZkbAvTsnyWDxT+MMjJ
GnEBVl4SULoMNMifiXPb/OBDR5rg/1CCe1VO29dYx+pBAzTTFfBjr6dL27vKK+imZkJsa0EFx7cs
7o7q2CyzuZ2lp0+wv4JGl1iqQsIK4Ji+5twXrt3kjSS72ejPim7HOJzXwcKwv1dO0pG5GuGuCuOg
Q0QQtDjaJOYP5Lr6LrCWI8YVlwUmL1GG+uQa13LiRGHzHZ6BcghItR8fVcbmZQCtD1S4ptnmFoPK
jECmGzIcZKhVE4ieDVR/2D0+iAMMVpKmHnFKdHrCB8SegEulGhLpK1ftrU6g1nLnQcz71MxRfM2t
DalItzh1NH4Wcw7dys3Vm6TfQ9DfyPBr7YtfhWoGBZouoT5p2bdwf2zOfUYkopcMsNnDS9EcVagM
oy08GRGDTvjhaXdeyV/funb3U2fFqRE408lpE7Yrha/hsN08lk49sQZejuwdc9iG195YNUhwk7TH
z1H8/M9mEMN0SIUg/sXgYllgP1qmyoC0qunk0NasIQ+EEoxIZtdOUcdPqstMutie2lPtobTr/GiD
R4NLm5E003UW3rRunJRpR2Jq28+Ly6yFOVtEVH+u2iiSDi6ud49+YLUAn32HHqrftn/TVK4Vw6ZH
PzKZh7SwKoZnc4+g9iuvXLrPMWDk8O/vsTHCA44rPNArXQES0DJHs2Vjtf527v81VcBMBZi/jqwf
ar39jdnoJSvVh5OlTbL2L0TZ/DPWv0Qw0mp9RpyBw1sWTV+tF0+jdyIXosTgx610SpsWgGtuoNic
Ok5WWzMeDL5WRlThaItYaSFoUaUf9KUrRzFz5JBGOXnstCNp16FgGY82lBIj7JbLJZUuAF6XU8eK
jAtL+xs7twHGC79VCLQj4WuaFHgHWrlN8arvYUW3TJ8PZYty11HVmLKsKZarT6MzsNFcA0dd5Yv2
1zjpi7YfAG9fNasJMHCWNbxi4mvQlRbbZVAznlRSTzTVcl+5z12ODAopKqGYDtnuW4fAEYhqowgA
bRaoE4rMuLOgahvok09SejYu66NxkAfUbUJDxZq0bjX9t858xEHcJ2Mf0OJHCDSsBS496UVKC1H5
Y1NxnTx0cidRtplmFNHnOYBECRMMxKqewbZt7iLwJKaxT4r+O6t7+2OItPOeJYyndTiRHRUSl5Wx
2vJYoPHzQBZAueExD7yFXuCT23hastLbQLZSNozv/4DVkebPfEk/0tvvmD4XoGV3H1OmD7yo/WfV
QU/Bmxg2IhPglUPu6M/XapCK6tqshXWMi/UV957R7uei9l4VqMtyMszW0CHrDOSXVAVAWqy1rwRR
mm4ubqaeJUJ6j5n9g95ZOcGdkXhwJPboy3ZCLq90SqxGkcJ01qMYOe9qQtrJNnNA9OmI/EDTtGS9
gOhwPFKJJIS6TM7x/tbcbumWhILIoC5GDScWEGX/UA5HAgP4Z3t80REXSalBrJy8YVqNT7vFomuI
6rt7K0fZMIDD8mY/0D72NYX7MvSLiHzlz79nUnF777CfwXoEUgDNL26yWFC3YlvbWvV48j7pO/D2
7VL2fm90BcCPnfNXr3QDJSPW55NHt5ePiLJ6+NWLC4bTtjCuy0ILChcDF/MyuE3DljIwH+qf6JF+
iG9f5gQOo1ot2ZE1fQ2MxMlBvkyuqDaqOGz32c0WV6xqrnOkbUH9AxaXQETHB3ebLoqihHWfH949
GUCV/nmzGbbzliAWM+uNNDZ0LsnRpRR9+2I1Km6sPouMwWgoHYUczSZ3M6yJE1aTDikSoklHege+
w53ZhJrvWYuKDZW5fvBHTkmCX1ioLAATAQu+gQvs0izfs+0WuD4axwm8kh3fjjTqO5WzrFeOfqu1
F+nD65HWgYFNryBAk6pPWdgKp8O2q6F1fS68WMjX3QSMdCY6Ox/W7/8AJ6vQDXaYlLmmDmBfU6Mw
tHWVcJy2OScwpIott5m4qMkJi1+H53utaeYddjJmDDXgNTiXwgGICHbqfOFjYIyWdIlos6/TOsw8
wi+VD3Emovx3OMMNXr9wCJJZhoqof0CmLZmD3pWuXoxMw8XV6bWzPBgq9uP23meExD9ZIR4hEgpS
V/qmHnjif4uYGejHktT1PV00VqrHrRAtPjheukmMHngLAZTPZ3BVoaJS2UjHHBfPzFEYd2At4YTS
9XNcZ55ePxDH+ckVs60rLeyD/p4CKlyUgEmWAm1fZhF9UiUJv8OGk2dqZySMAUrLQkR4LEKd1yY8
wpDvNHd0HqZq8VB5zib5zbvR9mwPsCJoGdgRfbULlLM75mIK/4OL7D2VAzQdfVY4r3WSLoYVYhXh
4KtCMKlaTv9ni0kjBrp4IGp26a+7Pkp12UAswT+r/XvNt0T38odSXumcHG94D8hFGSSH5D0QqAjt
/s+JGtF1orfeKxAcTOg4CWgB5+QuAfIJUZcD7wnjZZN3Zzp4Og8OShx2Qot/SzoxOIchjgBc+sjQ
Y0/lgdqxM/1bL7GB7SYsEbwIjj/qJJBf/L/hyaZPpF7Rlp24yP8whr8w8D/Sme80rQQwBftvCa9B
ku6+NLuTqYimTtjJHfXgpu7xSEI7O0uAgmzorTsgAylyul7gGxOpYkCUAhJ2nSGPMCxzXNtSXvfw
3glhceP5kaE0WDP6derqISICx33SCbm/mwLauLqsnPawT8TdRGlTweBGWhWbsG/wMWhIat38BV5X
lO/fI+JdyXFg4wHzA/mlfJwSWeXtPfsPxuS1AckpIDEcCOmoQV5DNqxzrrEWoZm9i65/kPPzcBOO
iiXY4M0UBmIGyViU9DVipaxjxHRcWekiIX63MQW+Pyo5+u5caXwlc9zOFasr7bOJJ8Bfb46IGS3z
YwQIWPks1eAbSZtCOeDcux+ciuqECdERKdfEYrYhFzVegQ6jKssCvhkMDgloiMzykWij+Nx5wNYj
/MX+Oq6Z+Mv01AoGt3PTqP+kqdI63N77UnkwsQPiZJtqm8jfVm7mREp60JU9TpqjxEW9YKikhZ1x
np0TqGWsD7SoJd0mYPaWoTSxt5AmyX1hwG8bHY51P8FcGjPq5nCwNi/AItFe8tebme9h5ZS4C6so
pAbWhsjdqoC7G46tyVp/mIYfvVJCPGGQz0xL9JnTbV9mHhSMVfEZpQ3ol3iWawaocfuTjcFyejqh
RtXq7vN7dVFQVZijytKKOBmKoR/W77yXjRbqIq6rtbNRLgHWozFnyWe4fj7ukwWJQ/futeFDocKq
85eZGPNflx5Daozgo/XiZ/WpdqKU8172NKmB50Ol+woQcgwNVIY+XtaXwvoLZdbj8unzWweYxuh3
n3FpNXhZy130c4W7Ly2HsSSp5SRNyGtIDk4iICKUIqRuS95oh2h9oJmE8bJ+4kgZsDWT+TbhnmIt
/p9fZBItGEhf7r4pAeEqarwc1ya1O9Zftmgmz0+6pmrvAqG6LXWfbtf3d6KkxjIxuL803snvg68D
PbxJdbugL0M3JeMEXcihoC8RhnisNEgOM4C70wnUNwH44j3pfK9iaJWHY99BprVlWoLTLnSQ7G9K
kWGy56nZGSt+f4eORbKF55hAnANZh6uHA4ihH4vy6trQVqY4qLtKT6EK+mOtHCd0f0FB+Br32U1r
5fXgrtH8A8JKR9LrL88WJh9ehRGfmp7S8I8mHZ6hHJsxf+cKwQr0T/1+ArTEtkIx0sfqv4stOzUS
NCsTDwzShafRn56n8JksjjptWkeVeOtkU5AdMPaIExPFztW+QNHzntJ9OxU55klXnLQJyTwJHW/q
KJyBVMM6aF+psdwTE6P6MT77PN6Aga7rgMGUK41tMYqMtVxsgW19GU7fCsNO3cwGZbjSV9DQHSs4
9MM9qhaOAKXdvK+KizN9Q1PX5bcoFzOkrdpF2Mv5JQgQDzZrqf15MkPnwVG3a86H4LgnjRKOWTpI
CnV3E6shFPRJriiV5Q8uhQ9sJP1tVd9aWc6rBsIcMyDbB+gJldfjS/wfJrI/m58YUgzqHZNXqFLt
SQcw4oD28P3yP6PUOilmBTA7yunsx9Dj3LOjw1m2RxOfl3jmg5dpcfEIqkxsI0Q2FkZ4vKiMBnSV
Vw5wQigqG9agEHgg4lxR4ij8aYsb+dTfoC8TGu7aUt4rUqaYSApLPeQQ6xjIYP4M+rDwPxqZuGKu
QmVqNloZEPLja8xv6rTE+Eaehlq6Oa69MJHgBYMbhvrJd9FzfQ8SaTrvmXlA45tnfB+4ya2e/f5L
A1mZMCee/N9GsWaN+i4+A2m/VfSyd/RYwComQrNkzdQzdncGFjCLwoSkDt4XNBCagGfX//03o0S1
OR4l5gOrHpYe3cuBlaWAAqVbSGcN6Tof5PxmgHXT7JU38XEm6aNPm9H+JW6tL3oOCHt7jeuofxf8
C5KzTfFGwUqcI6l81/UTjKOLD+GjvPHCOlboEuIBoER46Rgbut+CqCVKxWWGzR4PW4KXZPULebVq
eqOX1MQwSDcuIhe1lkDZYHGomJmKZVhxh3syX24VCxsmja7KC2VNHcHcfsinE+45DLXtKalu2FQ8
d8VsJUju1vzS+5PMw9bj+gHNAgu+9+nvKLnijACWxopd1fTcMjZ1/DafcmVw7i+O5A+kue3DgX6f
bdQe8XPMNQgJEtU3f9rEIKJ+9rtD1ry7NRd9I88GA+MGYVDMAlAuPclnhPO+/0c8e4852JSzFUsM
D9pmwykUayOb5H/mq34YWoYlSM0sPi+Qm0GIS4iRqPchZSIakDmKI0C5a5US8A/qxKKdDyGEVZ58
p3ndF0VxAe2pdjeQ1UkIRIuh2pl9+Ub9zfPAjhLbMi8kBoGynnPc1wkbD8pFJsbAJc4TpccwOqVh
/g2zLaW2DDVkPvgkdv36PS1TNw6XhCMKuKBvwEbeaN3H/oGgYMQhLtboqZA2pTKoxYrY49NXjORS
EnDxg8WTOgIo6FfjOE9DlgiN1rIa6V7GwjNV3v5HlLCKeyu1/9hBSpMXfvRZ+SypHTJ792rqjNnN
dyCLemHQ3F1WzM1X7szELyVQuOsU5SzmHGPxgk7NH5SAhjCwu17PxMlJlu3iGkcXSulQox+86IKM
egwrVIIYO9zRL/rSGdGwM2dCWNtihN0Oo/W+Zdw2lcD/GfvGWwzwkdFQ37YsjWTmklCzozDpybtD
9XJfRChBuFXNIatqV+Tw/k4XK/VowHPE6Mh5GdcuoDv0SOvQTpN2dK3VGiAdvcGouXiL4UXoiinW
odueFlb0D+Hya1UB3NBob4U5lH9bAPTGIuhcDlS9A9NNjtXtmr97KGuzXThNkpi6TNTbia6NAyGs
6awm9n2tuJtPvA7WV5spbIYRZl3mCL8G1j/e5YHTaKqW++ovpKxGzuLl8nc2oNRuEVn+JRabGgLZ
iv5ZXWlSFO8YrJSFfE2s6yl2qk7cHiytSWd5vRMA71tzCdH8DrxR9fEnSpRDbqeG3/LkZ8ZolT+i
NstfHwXrrLLL/XezSROSXrOiPQ0XsQJHLt7NWgDqz8RsGzepbyW+keTqMD7ZzXXf40/nOVmBbGGO
hURZE1/dyY4eStqKfikvGWVemyEE+yWrfSa5MSDOUbqovyAxLjA4nwGwsvES7C2xEjs52xAD7dFE
VgUtKvLZPEXimiBk8GT9fT6/GYhxLBewiFb+eIJLguEd8OiIv62141It3jppiZ6RaoAHkADf36Oj
wNWL8bF7YztIJKPNoLhbksFxSMeDo+kJ8n40lrisU7+tlOke4CWGzwfwCAE6qH7CEpb/HZWjRT1+
llBA+SdKlhpDXpL2FNzpQRQm5hMei+CORJFdwb5fjvAUDXN9lnWESIGSXuKUj+86SjfbCEit4LR7
P5Ymm1kRtdguPW7vvFguvO6OMVezIntctNtZHknJTW0Ovd5Sfcyt0JnrkIje5C9S+fBSM1LQ4jM4
Zszo5gaU8Bm3T0RSYYJp8LViDvOPze4PaWfXQLyQvQRml5AhdcpcN7e7g6/ywtUCdVnxvnx0Z1CP
fhyg5g2882eIrg27Wesi32rQnPyj7y88ubicijsaxn24LIszp20OnrXI2OL+QrIdZvx3DoX7CsFx
dR607UAtdbbghN2HK0q3b+p2Z4RAK6MXYLeyy+1PLlHbRqumC0pkzqxktJzNpHghDzLMiM49c40V
aAZOwnhsX1pn3LASLwPUPFqSnIWcXGicJrXawp5+7uqlB9XmADUU6/0H2MwBix+YkM4rzjoXU/4x
/ef5WkjoBFbppfTDcDd47dKZIC4XWDffqPcNbMoj1Tdzc68CXAnvL2EVQCB19G1yqHAX+HiiEmw9
3MK4FRdt70Ucft7VIMZFFC106oOFoD5if0ckk21xJC7AOULQhNgLDc5+3/b73ArfInaHrTI2nTN3
TWFPk4w8sd+vCkLCG4XWeUnqPUNI/QM87y1ABDBmKaTnhc2QibcBiJrXi8JOn8CzNYVMXm2kRUkp
TuifuhKpFtEZ5ErUJcRgWYqOpKeHRxF11Ca2gW368V6k7jL6y7jKtGZKJWGpndXCABGeRMRHJAll
50qTqu1gKV1tNU3kGXWgCvlq622Rwl5Mtx1xvtWgtFBbtRsTxVmtkJ73iG8fcOLSX7m90EYfVEcr
ALQutxzWPfKTrXSiLga8s9Gx/obiujpDXdmFJslLk4VA0b7parDPR4W+SFBTMpBjO1dE3saO3Hgw
6JHe0UUOQNEtCx35bJLWMRLUFAVbaAzUSPdMzMPdVpJuBf+xN/XUKxggJJrlhGb3OgHlUStz+nYJ
1loe5pM7whMJtG3iVZz3s1VjPp6y76jvEOWdcqzxGV1gYo7+Spn2ztG+YdoHEBwvwGO60kvVY0mW
U7W09tvAkH85t/1s+SbkhlaccwAOY1X91rYfwJSNRFQCSoImEUBl0o7/E8zhv8oJ7ZOMcjqyI+tE
t1eSkYKw8b7MH2qsPoWLvWJUc89I5rZFKPf1V54WyoXK408Wydke9oE2dc2wPvFPtThApYNOl4/Y
ITxfs2kjmrSo+xp/PiM3X9C90wKc6Uqv4fpAxiROXrbKCfntiBPxiANDFw4HhK87ZjSKkSRUVR7K
ozuRJ+EH8AuU9+dMf7KpB4TD7ZmER2A5ENKqVZf3RTYC4jTXJnM8WrhjYxIBTKXw89AJSwkII/Eb
9lK4l/RTEnRMcOMWaLbeKTPQuLwFXGVA2KVDJkGyBZh5AlcNLsGJCsDp2oWWoQ7w2uhFdOpYrhlt
nBQ8yzIzCUIVQtfWUpFE2o7+oKM7q+CkKI7nbE5/LKp81k+g23rpGuXO/7jNoyaJ4nCzpsu/1Dhc
CXO2DMyX2rTM+dqRdxVOMz/vawU/06LD2TeVr752ckgklmB6Cm3FYGisQRhlV0lpGRZnhG6H45QW
1ml5a7DRgT0H182vwy8vHnEmOjtL9bl1hxOUhg0D+FDhH0E/ZczxqZGQhOLTe+L31dPjuwkOBshA
fOKOsjyVy+IiJmkdi+i8rTlYJQFE6zljpJKvQS9BC6/OkFSIOMsSJv5CeDp0cqU6GNETZBALlzny
sPyvYN6OMvHEvdKerJSN36uwX8u1Nn4JW0c8r2OlkhPAV+9wU3yE5thMQKG5AaVStDJDzQf3+Cu+
D7KcEeJQc9/Dsd/njl+x06s6ImtnbtVyKvKZIOTrT49YuUImHoZzutrzaNhb/vb7POP2tvxFc6YG
Tmk3wBB72G9dfrUKd1RVVkrteDAvvvRlEubIMHaAhL9Zn55CmhaKj6TNl0tXY1XzCOmOwgeyObA3
07tLAOa4fsPkTRwsUM2EfQ+3XlLwJEgFAWg0Bi7nRkRa60T8m1DS2uycn0xSOFRwKbN7VTiDA0Ut
h3FPLepMNu/qtwvb/qDQgCbNbX+9G7jFav6w3W0VGc//2MUqCRI+q+aXYeB33atz5fQeb8ro1dzd
nwDsTZiBaG5fjBU15IExoObjZmx5TAldDmXsnfYV9PsnInlzpAznGnX69MaHHdnZOsm1JZCsMdzX
n4e3atadf6dKh7RH54LKyZUtfkBqg4ga4vM63iXJ8463lzOpXnx025OvkAXFb/1b9IpZ/pN9mJGg
OFVCYtaoxfokjn9nzAqv6YQvDFADBbVEFvE6F5PaaeXCZs+CKSP4Qx6CWqkUAftuktU+M9gsHPOa
y4LVTdKAswJux2DEqw1OEL/hGNSF8xtyaE8O/+yuIzU9YS11GNr7mh9SF28dxzwPCi7CK71r76cn
07ygR3z/OLJXRmGv2HsEaVWYrxvs3IxTkZwC223kStIKJuGFGDzXznToVnMp3GSNqc+EDDVyUM5y
lV8YC2bwADIoHoz1QzYS4LlCFjZPwL1Azy55b8TD9q6Fy8LpmQHuwMI3xlmI3nauAlOmTG4xSP3q
0aKonlC3kM+kbD5bKWtqOzen/l0cCUPFdav4uUghOnaTg3aVF/Dc2Cu2KPacHkU6OR+yshOzE6YH
95IWSH8FcQz2VmOGEvYS/7iftiYYS+VejwHrnYnvJwWprd54wh0KPs+WAhEgttoU23pg6nsfhzGI
PcRz5qEakH3N53KT4QvUvPc56QzZi1IAhNe0XHroGFHwso8PDu4dehfoKZ9jBdTke27SAODCwpyK
Q2ELBnN/SZX8TXv9zfm3J/mMjqyPcE//NzIXKd5ATZDHRdzNX50MvgpOOOpoVCOwpSQN9qKtlYLK
0i2h/tg4w03eEOBxUXSsqWTbqYEzXGa+5n1QahEm54lGcB1pkzN3qFeF+AAIceA/l3qg3qzLVBg4
B0mx/l7FKkEy8poWRFRKfq713+MvTBtPCDbEOMCnx2ltsLczDiwdvUXR7g7XLcLyxBkMX93U4JIy
PC/PscDTAxFGo8GhJ4npwyyPhYsNFDJvJEDn9UlYJ3GvetLxnBHo6f6E/xadZQI6JSzolhxV4+8K
2Afk7Mq6srG/R55KagGW8ll6LjshCC+1u/krBBC4a5HgBwwQGycl62r192T1ad5o1l8/OHprIy9I
TPMWXtYjmZKJ2Jk3xvKnsQEcNwpozDAhtuKbV+rvGofVodpVdCiaSYq4xCP7faibsx2GSOHNAuTJ
F3vsqG22Px4aq+UuiDR5dxG8+9PCYHRRRLYYL+wZVtBTpQvZUuyCngixp0cnQxiFR95cx0m70rH9
nWwxR0HCOG0sopSuj069BSJaGBMoAFzbOwyriYIU1P8wSI6+WRiN5PC0yysbgm2EM/XU7Q9Xi1yW
b+6ukZrEK2kybFJnbaj8VhoqcsRE6SDk+UkBBHPQdCZpl+QzWtK4fdbi2lFGMzIy2/LhGzffNBOL
cxmnYrtEVBrdJe5dDqL7tjZQre0=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity FIFO_SC_HS_Top is
port(
  Data :  in std_logic_vector(7 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(7 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end FIFO_SC_HS_Top;
architecture beh of FIFO_SC_HS_Top is
  signal Clk_d : std_logic ;
  signal WrEn_d : std_logic ;
  signal RdEn_d : std_logic ;
  signal Reset_d : std_logic ;
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal Full_d : std_logic ;
  signal Empty_d : std_logic ;
  signal Data_d : std_logic_vector(7 downto 0);
  signal Q_d : std_logic_vector(7 downto 0);
component \~fifo_sc_hs.FIFO_SC_HS_Top\
port(
  Clk_d: in std_logic;
  Reset_d: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn_d: in std_logic;
  RdEn_d: in std_logic;
  Data_d : in std_logic_vector(7 downto 0);
  Full_d: out std_logic;
  Empty_d: out std_logic;
  Q_d : out std_logic_vector(7 downto 0));
end component;
begin
Data_0_ibuf: IBUF
port map (
  O => Data_d(0),
  I => Data(0));
Data_1_ibuf: IBUF
port map (
  O => Data_d(1),
  I => Data(1));
Data_2_ibuf: IBUF
port map (
  O => Data_d(2),
  I => Data(2));
Data_3_ibuf: IBUF
port map (
  O => Data_d(3),
  I => Data(3));
Data_4_ibuf: IBUF
port map (
  O => Data_d(4),
  I => Data(4));
Data_5_ibuf: IBUF
port map (
  O => Data_d(5),
  I => Data(5));
Data_6_ibuf: IBUF
port map (
  O => Data_d(6),
  I => Data(6));
Data_7_ibuf: IBUF
port map (
  O => Data_d(7),
  I => Data(7));
Clk_ibuf: IBUF
port map (
  O => Clk_d,
  I => Clk);
WrEn_ibuf: IBUF
port map (
  O => WrEn_d,
  I => WrEn);
RdEn_ibuf: IBUF
port map (
  O => RdEn_d,
  I => RdEn);
Reset_ibuf: IBUF
port map (
  O => Reset_d,
  I => Reset);
Q_0_obuf: OBUF
port map (
  O => Q(0),
  I => Q_d(0));
Q_1_obuf: OBUF
port map (
  O => Q(1),
  I => Q_d(1));
Q_2_obuf: OBUF
port map (
  O => Q(2),
  I => Q_d(2));
Q_3_obuf: OBUF
port map (
  O => Q(3),
  I => Q_d(3));
Q_4_obuf: OBUF
port map (
  O => Q(4),
  I => Q_d(4));
Q_5_obuf: OBUF
port map (
  O => Q(5),
  I => Q_d(5));
Q_6_obuf: OBUF
port map (
  O => Q(6),
  I => Q_d(6));
Q_7_obuf: OBUF
port map (
  O => Q(7),
  I => Q_d(7));
Empty_obuf: OBUF
port map (
  O => Empty,
  I => Empty_d);
Full_obuf: OBUF
port map (
  O => Full,
  I => Full_d);
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.FIFO_SC_HS_Top\
port map(
  Clk_d => Clk_d,
  Reset_d => Reset_d,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn_d => WrEn_d,
  RdEn_d => RdEn_d,
  Data_d(7 downto 0) => Data_d(7 downto 0),
  Full_d => Full_d,
  Empty_d => Empty_d,
  Q_d(7 downto 0) => Q_d(7 downto 0));
end beh;
