
module sid_tables
#(
	parameter MULTI_FILTERS   = 1
)
(
	input             clock,
	input             mode,

	// waves
	input      [11:0] acc_t,
	output reg  [7:0] _st_out,
	output reg  [7:0] p_t_out,
	output reg  [7:0] ps__out,
	output reg  [7:0] pst_out,

	// filter
	input       [1:0] cfg,
	input      [10:0] Fc,
	input      [12:0] Fc_offset,
	output     [15:0] F0,
	input             ld_clk,
	input      [11:0] ld_addr,
	input      [15:0] ld_data,
	input             ld_wr
);

// P + T
always_ff @(posedge clock) begin
	p_t_out <= mode ? wave8580_p_t[acc_t[10:0]] : wave6581_p_t[acc_t[10:0]];
end

// P + S
always_ff @(posedge clock) begin
	ps__out <= mode ? wave8580_ps_[acc_t] : wave6581_ps_[acc_t[10:0]];
end

// S + T
always_ff @(posedge clock) begin
	_st_out <= mode ? {
		((acc_t & 'he7e) == 'he7e) | ((acc_t & 'he80) == 'he80) | ((acc_t & 'hf00) == 'hf00) | ((acc_t & 'he7d) == 'he7d),
		((acc_t & 'h7f8) == 'h7f8) | ((acc_t & 'hf00) == 'hf00),
		((acc_t & 'h7e0) == 'h7e0) | ((acc_t & 'hf0f) == 'hf0f) | ((acc_t & 'hf1b) == 'hf1b) | ((acc_t & 'hbfe) == 'hbfe) | ((acc_t & 'hf1e) == 'hf1e) | ((acc_t & 'hf40) == 'hf40) | ((acc_t & 'hf30) == 'hf30) | ((acc_t & 'hf29) == 'hf29) | ((acc_t & 'hf26) == 'hf26) | ((acc_t & 'hf80) == 'hf80),
		((acc_t & 'h7e0) == 'h7e0) | ((acc_t & 'h3f0) == 'h3f0) | ((acc_t & 'hdfe) == 'hdfe) | ((acc_t & 'h5ff) == 'h5ff) | ((acc_t & 'hf80) == 'hf80),
		((acc_t & 'h7e0) == 'h7e0) | ((acc_t & 'h3f0) == 'h3f0) | ((acc_t & 'hfc0) == 'hfc0) | ((acc_t & 'h1f8) == 'h1f8) | ((acc_t & 'heff) == 'heff),
		((acc_t & 'h0fc) == 'h0fc) | ((acc_t & 'h1f8) == 'h1f8) | ((acc_t & 'h3f0) == 'h3f0) | ((acc_t & 'hfe0) == 'hfe0),
		((acc_t & 'h07e) == 'h07e) | ((acc_t & 'hff0) == 'hff0) | ((acc_t & 'h7f7) == 'h7f7) | ((acc_t & 'h1f8) == 'h1f8) | ((acc_t & 'h0fc) == 'h0fc),
		((acc_t & 'hdbf) == 'hdbf) | ((acc_t & 'h0fc) == 'h0fc) | ((acc_t & 'h3fa) == 'h3fa) | ((acc_t & 'h7f8) == 'h7f8) | ((acc_t & 'h3bf) == 'h3bf) | ((acc_t & 'h07e) == 'h07e)
	} : {
		1'b0,
		((acc_t & 'h7fc) == 'h7fc),
		((acc_t & 'h7e0) == 'h7e0) | ((acc_t & 'h3fe) == 'h3fe),
		((acc_t & 'h7e0) == 'h7e0) | ((acc_t & 'h5ff) == 'h5ff) | ((acc_t & 'h3f0) == 'h3f0),
		((acc_t & 'h7e0) == 'h7e0) | ((acc_t & 'h1f8) == 'h1f8) | ((acc_t & 'h3f0) == 'h3f0),
		((acc_t & 'h0fc) == 'h0fc) | ((acc_t & 'h1f8) == 'h1f8) | ((acc_t & 'h3f0) == 'h3f0),
		((acc_t & 'h07e) == 'h07e) | ((acc_t & 'h1f8) == 'h1f8) | ((acc_t & 'h0fc) == 'h0fc),
		((acc_t & 'h13f) == 'h13f) | ((acc_t & 'h07e) == 'h07e) | ((acc_t & 'h7fa) == 'h7fa) | ((acc_t & 'h0bf) == 'h0bf) | ((acc_t & 'h0fc) == 'h0fc)
	};
end

// P + S + T
always_ff @(posedge clock) begin
	pst_out <= mode ? {
		((acc_t & 'he89) == 'he89) | ((acc_t & 'he3e) == 'he3e) | ((acc_t & 'hec0) == 'hec0) | ((acc_t & 'he8a) == 'he8a) | ((acc_t & 'hdf7) == 'hdf7) | ((acc_t & 'hdf8) == 'hdf8) | ((acc_t & 'he85) == 'he85) | ((acc_t & 'he6a) == 'he6a) | ((acc_t & 'he90) == 'he90) | ((acc_t & 'he83) == 'he83) | ((acc_t & 'he67) == 'he67) | ((acc_t & 'hea0) == 'hea0) | ((acc_t & 'hf00) == 'hf00) | ((acc_t & 'he5e) == 'he5e) | ((acc_t & 'he70) == 'he70) | ((acc_t & 'he6c) == 'he6c),
		((acc_t & 'heee) == 'heee) | ((acc_t & 'h7ef) == 'h7ef) | ((acc_t & 'h7f2) == 'h7f2) | ((acc_t & 'h7f4) == 'h7f4) | ((acc_t & 'hef0) == 'hef0) | ((acc_t & 'h7f8) == 'h7f8) | ((acc_t & 'hf00) == 'hf00) | ((acc_t & 'h7f1) == 'h7f1),
		((acc_t & 'hf78) == 'hf78) | ((acc_t & 'h7f0) == 'h7f0) | ((acc_t & 'h7ee) == 'h7ee) | ((acc_t & 'hf74) == 'hf74) | ((acc_t & 'hf6f) == 'hf6f) | ((acc_t & 'hf80) == 'hf80) | ((acc_t & 'hbff) == 'hbff),
		((acc_t & 'hdff) == 'hdff) | ((acc_t & 'hbfe) == 'hbfe) | ((acc_t & 'h7ef) == 'h7ef) | ((acc_t & 'h7f2) == 'h7f2) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'h7f4) == 'h7f4) | ((acc_t & 'hfc0) == 'hfc0) | ((acc_t & 'hfb8) == 'hfb8) | ((acc_t & 'h7f8) == 'h7f8) | ((acc_t & 'hfb6) == 'hfb6),
		((acc_t & 'hbfe) == 'hbfe) | ((acc_t & 'hfdc) == 'hfdc) | ((acc_t & 'hdfe) == 'hdfe) | ((acc_t & 'h7f7) == 'h7f7) | ((acc_t & 'hfda) == 'hfda) | ((acc_t & 'hbfd) == 'hbfd) | ((acc_t & 'h7f8) == 'h7f8) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'hfe0) == 'hfe0) | ((acc_t & 'heff) == 'heff),
		((acc_t & 'hfeb) == 'hfeb) | ((acc_t & 'h7fa) == 'h7fa) | ((acc_t & 'hbfe) == 'hbfe) | ((acc_t & 'hdfe) == 'hdfe) | ((acc_t & 'hff0) == 'hff0) | ((acc_t & 'h7fc) == 'h7fc) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'hfec) == 'hfec) | ((acc_t & 'heff) == 'heff),
		((acc_t & 'hff6) == 'hff6) | ((acc_t & 'hdff) == 'hdff) | ((acc_t & 'hf7f) == 'hf7f) | ((acc_t & 'hbfe) == 'hbfe) | ((acc_t & 'h7fc) == 'h7fc) | ((acc_t & 'hff5) == 'hff5) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'hff8) == 'hff8) | ((acc_t & 'heff) == 'heff),
		((acc_t & 'hdff) == 'hdff) | ((acc_t & 'hf7f) == 'hf7f) | ((acc_t & 'hffa) == 'hffa) | ((acc_t & 'h7fe) == 'h7fe) | ((acc_t & 'hff9) == 'hff9) | ((acc_t & 'hffc) == 'hffc) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'heff) == 'heff)
	} : {
		1'b0,
		((acc_t & 'h7fc) == 'h7fc) | ((acc_t & 'h7fb) == 'h7fb),
		((acc_t & 'h7ef) == 'h7ef) | ((acc_t & 'h7f7) == 'h7f7) | ((acc_t & 'h7fc) == 'h7fc) | ((acc_t & 'h7fb) == 'h7fb) | ((acc_t & 'h3ff) == 'h3ff),
		((acc_t & 'h7fc) == 'h7fc) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'h7f7) == 'h7f7) | ((acc_t & 'h7fb) == 'h7fb),
		((acc_t & 'h7fc) == 'h7fc) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'h7fb) == 'h7fb),
		((acc_t & 'h7fd) == 'h7fd) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'h7fe) == 'h7fe),
		((acc_t & 'h7fd) == 'h7fd) | ((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'h7fe) == 'h7fe),
		((acc_t & 'h3ff) == 'h3ff) | ((acc_t & 'h7fe) == 'h7fe)
	};
end


wire [7:0] wave6581_p_t[0:2047] = 
'{
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h20, 'h38, 'h3f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h40, 'h40, 'h5f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h00, 'h00, 'h60, 'h00, 'h60, 'h60, 'h6f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60, 'h00, 'h00, 'h00, 'h60, 'h00, 'h60, 'h70, 'h77,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60, 'h00, 'h00, 'h00, 'h70, 'h40, 'h70, 'h70, 'h7b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h70, 'h00, 'h40, 'h40, 'h70, 'h60, 'h70, 'h78, 'h7d,
	'h00, 'h40, 'h60, 'h78, 'h60, 'h78, 'h78, 'h7e, 'h70, 'h7c, 'h7c, 'h7f, 'h7e, 'h7f, 'h7f, 'h7f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h9f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'h80, 'h80, 'ha0, 'ha0, 'haf,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'ha0, 'h00, 'h80, 'h80, 'ha0, 'h80, 'ha0, 'hb0, 'hb7,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'ha0,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'ha0, 'h00, 'h80, 'h80, 'ha0, 'h80, 'hb0, 'hb0, 'hbb,
	'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'hb0, 'h80, 'h80, 'h80, 'hb0, 'h80, 'hb0, 'hb8, 'hbd,
	'h80, 'h80, 'h80, 'hb8, 'ha0, 'hb8, 'hb8, 'hbe, 'ha0, 'hb8, 'hbc, 'hbf, 'hbe, 'hbf, 'hbf, 'hbf,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'hc0,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h80, 'hc0,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'hc0,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'hc0, 'h00, 'h80, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hcf,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'hc0,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'hc0,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'hc0, 'hc0, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd0, 'hd7,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'hc0, 'hc0,
	'h00, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'hc0, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hd0, 'hd0, 'hdb,
	'h00, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'hd0, 'h80, 'hc0, 'hc0, 'hd0, 'hc0, 'hd0, 'hd8, 'hdd,
	'hc0, 'hc0, 'hc0, 'hd0, 'hc0, 'hd8, 'hd8, 'hde, 'hc0, 'hd8, 'hdc, 'hdf, 'hdc, 'hdf, 'hdf, 'hdf,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h80, 'hc0, 'hc0, 'he0,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'he0,
	'h00, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'he0, 'h80, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'he7,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'hc0, 'h00, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'he0,
	'h00, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'he0, 'hc0, 'hc0, 'hc0, 'he0, 'he0, 'he0, 'he0, 'heb,
	'h80, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'hed,
	'hc0, 'he0, 'he0, 'he0, 'he0, 'he8, 'he8, 'hee, 'he0, 'he8, 'hec, 'hef, 'hec, 'hef, 'hef, 'hef,
	'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'hc0, 'h80, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hf0,
	'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'he0, 'hf0, 'hc0, 'he0, 'he0, 'hf0, 'he0, 'hf0, 'hf0, 'hf3,
	'h80, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'hf0, 'hc0, 'he0, 'he0, 'hf0, 'he0, 'hf0, 'hf0, 'hf5,
	'he0, 'he0, 'he0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf6, 'hf0, 'hf0, 'hf4, 'hf7, 'hf4, 'hf7, 'hf7, 'hf7,
	'hc0, 'hc0, 'hc0, 'he0, 'he0, 'he0, 'he0, 'hf0, 'he0, 'he0, 'he0, 'hf8, 'hf0, 'hf8, 'hf8, 'hf9,
	'he0, 'hf0, 'hf0, 'hf8, 'hf0, 'hf8, 'hf8, 'hfa, 'hf0, 'hf8, 'hf8, 'hfb, 'hf8, 'hfb, 'hfb, 'hfb,
	'he0, 'hf0, 'hf0, 'hf8, 'hf0, 'hf8, 'hfc, 'hfc, 'hf8, 'hfc, 'hfc, 'hfd, 'hfc, 'hfd, 'hfd, 'hfd,
	'hf8, 'hfc, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff
};


wire [7:0] wave6581_ps_[0:2047] = 
'{
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h07,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h02, 'h1f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h2f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h37,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3d,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3e,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h30, 'h3f, 'h00, 'h30, 'h38, 'h3f, 'h3e, 'h3f, 'h3f, 'h3f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h4f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h57,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h5b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h5d,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h5e,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h5f, 'h00, 'h40, 'h40, 'h5f, 'h5c, 'h5f, 'h5f, 'h5f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h67,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h6b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h40, 'h6d,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h00, 'h00, 'h40, 'h00, 'h40, 'h40, 'h6e,
	'h00, 'h00, 'h00, 'h40, 'h00, 'h60, 'h60, 'h6f, 'h00, 'h60, 'h60, 'h6f, 'h60, 'h6f, 'h6f, 'h6f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h00, 'h00, 'h40, 'h00, 'h40, 'h60, 'h73,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h00, 'h00, 'h40, 'h00, 'h60, 'h60, 'h75,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60, 'h00, 'h00, 'h00, 'h60, 'h00, 'h60, 'h60, 'h76,
	'h00, 'h00, 'h00, 'h60, 'h00, 'h60, 'h60, 'h77, 'h00, 'h70, 'h70, 'h77, 'h70, 'h77, 'h77, 'h77,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60, 'h00, 'h00, 'h00, 'h60, 'h00, 'h60, 'h60, 'h79,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h60, 'h00, 'h00, 'h00, 'h60, 'h00, 'h70, 'h70, 'h7a,
	'h00, 'h00, 'h00, 'h70, 'h00, 'h70, 'h70, 'h7b, 'h40, 'h70, 'h70, 'h7b, 'h78, 'h7b, 'h7b, 'h7b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h70, 'h00, 'h00, 'h00, 'h70, 'h00, 'h70, 'h70, 'h7c,
	'h00, 'h00, 'h00, 'h70, 'h40, 'h70, 'h70, 'h7d, 'h40, 'h70, 'h78, 'h7d, 'h78, 'h7d, 'h7d, 'h7d,
	'h00, 'h40, 'h40, 'h78, 'h60, 'h78, 'h78, 'h7e, 'h60, 'h78, 'h78, 'h7e, 'h7c, 'h7e, 'h7e, 'h7e,
	'h70, 'h7c, 'h7c, 'h7f, 'h7e, 'h7f, 'h7f, 'h7f, 'h7e, 'h7f, 'h7f, 'h7f, 'h7f, 'h7f, 'h7f, 'h7f
};


wire [7:0] wave8580_p_t[0:2047] =
'{
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h07,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h1c, 'h00, 'h3c, 'h3f, 'h3f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h0c, 'h5e, 'h5f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h00, 'h00, 'h40, 'h40, 'h60, 'h60, 'h6f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h40,
	'h00, 'h00, 'h00, 'h40, 'h40, 'h40, 'h40, 'h60, 'h40, 'h40, 'h60, 'h60, 'h60, 'h60, 'h70, 'h77,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h40, 'h40, 'h40, 'h40, 'h40, 'h40, 'h40, 'h60, 'h60, 'h60,
	'h40, 'h40, 'h40, 'h60, 'h60, 'h60, 'h60, 'h70, 'h60, 'h60, 'h60, 'h70, 'h70, 'h70, 'h78, 'h7b,
	'h60, 'h60, 'h60, 'h70, 'h60, 'h70, 'h70, 'h70, 'h70, 'h70, 'h70, 'h78, 'h78, 'h78, 'h78, 'h7c,
	'h78, 'h78, 'h78, 'h7c, 'h78, 'h7c, 'h7c, 'h7e, 'h7c, 'h7e, 'h7e, 'h7f, 'h7f, 'h7f, 'h7f, 'h7f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h8e, 'h9f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'h80,
	'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'haf,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'ha0, 'ha0, 'ha0, 'ha0, 'hb7,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'ha0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'ha0, 'ha0, 'ha0, 'ha0, 'ha0, 'hb0, 'ha0, 'hb0, 'hb0, 'hbb,
	'ha0, 'ha0, 'ha0, 'ha0, 'ha0, 'ha0, 'hb0, 'hb0, 'ha0, 'hb0, 'hb0, 'hb8, 'hb0, 'hb8, 'hb8, 'hbc,
	'hb0, 'hb8, 'hb8, 'hb8, 'hb8, 'hbc, 'hbc, 'hbe, 'hbc, 'hbc, 'hbe, 'hbf, 'hbe, 'hbf, 'hbf, 'hbf,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'hc0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'h80, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'h80, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hcf,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'hc0, 'hc0, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd7,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd0, 'hd0, 'hd9,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd0, 'hc0, 'hd0, 'hd0, 'hd0, 'hd0, 'hd8, 'hd8, 'hdc,
	'hd0, 'hd0, 'hd8, 'hd8, 'hd8, 'hdc, 'hdc, 'hde, 'hdc, 'hdc, 'hde, 'hdf, 'hde, 'hdf, 'hdf, 'hdf,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'he0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'hc0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he7,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he8,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he8, 'hec,
	'he0, 'he0, 'he0, 'he8, 'he8, 'he8, 'hec, 'hee, 'hec, 'hec, 'hec, 'hee, 'hee, 'hef, 'hef, 'hef,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'hf0, 'hf0, 'hf0,
	'he0, 'he0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0,
	'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf4,
	'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf4, 'hf0, 'hf4, 'hf4, 'hf6, 'hf6, 'hf7, 'hf7, 'hf7,
	'hf0, 'hf0, 'hf0, 'hf8, 'hf0, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8,
	'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hfa, 'hfa, 'hfb, 'hfb, 'hfb,
	'hf8, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfd, 'hfd, 'hfd,
	'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff
};


wire [7:0] wave8580_ps_[0:4095] =
'{
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h0f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h07,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h07, 'h07, 'h1f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01, 'h0f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h17,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3d,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3e,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h3f, 'h00, 'h0c, 'h1c, 'h3f, 'h1e, 'h3f, 'h3f, 'h3f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h0f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h07,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h0b,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h0a,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h5e,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h5f, 'h00, 'h00, 'h00, 'h5f, 'h0c, 'h5f, 'h5f, 'h5f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h47,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h43,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h65,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h6e,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h6f, 'h00, 'h40, 'h40, 'h6f, 'h40, 'h6f, 'h6f, 'h6f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h63,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h61,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h00, 'h00, 'h00, 'h40, 'h00, 'h40, 'h40, 'h70,
	'h00, 'h00, 'h40, 'h40, 'h40, 'h40, 'h40, 'h70, 'h40, 'h60, 'h60, 'h77, 'h60, 'h77, 'h77, 'h77,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h40, 'h60, 'h00, 'h40, 'h40, 'h60, 'h40, 'h60, 'h60, 'h79,
	'h00, 'h40, 'h40, 'h40, 'h40, 'h40, 'h40, 'h60, 'h40, 'h40, 'h40, 'h60, 'h60, 'h60, 'h60, 'h78,
	'h40, 'h60, 'h60, 'h60, 'h60, 'h60, 'h60, 'h78, 'h60, 'h70, 'h70, 'h78, 'h70, 'h79, 'h7b, 'h7b,
	'h60, 'h60, 'h60, 'h60, 'h60, 'h60, 'h60, 'h70, 'h60, 'h60, 'h60, 'h70, 'h60, 'h70, 'h70, 'h7c,
	'h60, 'h70, 'h70, 'h70, 'h70, 'h70, 'h70, 'h7c, 'h70, 'h78, 'h78, 'h7c, 'h78, 'h7c, 'h7c, 'h7d,
	'h70, 'h78, 'h78, 'h78, 'h78, 'h78, 'h78, 'h7c, 'h78, 'h7c, 'h7c, 'h7e, 'h7c, 'h7e, 'h7e, 'h7e,
	'h7c, 'h7c, 'h7c, 'h7e, 'h7e, 'h7f, 'h7f, 'h7f, 'h7e, 'h7f, 'h7f, 'h7f, 'h7f, 'h7f, 'h7f, 'hff,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h03,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h8f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h87,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h83,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h8d,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'h8e,
	'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h8f, 'h80, 'h80, 'h80, 'h9f, 'h80, 'h9f, 'h9f, 'h9f,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h01,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h80, 'h80, 'h87,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h83,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h81,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h84,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h87, 'h80, 'h80, 'h80, 'h87, 'h80, 'h8f, 'haf, 'haf,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h80, 'h80, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h83,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h81,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'ha0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'ha0, 'h80, 'h80, 'h80, 'ha0, 'h80, 'ha3, 'hb7, 'hb7,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hb1,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hb0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hb0, 'h80, 'ha0, 'ha0, 'hb0, 'ha0, 'hb8, 'hb9, 'hbb,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'ha0, 'h80, 'h80, 'h80, 'ha0, 'h80, 'ha0, 'ha0, 'hb8,
	'h80, 'ha0, 'ha0, 'ha0, 'ha0, 'ha0, 'ha0, 'hb8, 'ha0, 'hb0, 'hb0, 'hb8, 'hb0, 'hbc, 'hbc, 'hbd,
	'ha0, 'hb0, 'hb0, 'hb0, 'hb0, 'hb8, 'hb8, 'hbc, 'hb0, 'hb8, 'hb8, 'hbc, 'hb8, 'hbc, 'hbe, 'hbe,
	'hb8, 'hbc, 'hbc, 'hbe, 'hbc, 'hbe, 'hbe, 'hbf, 'hbe, 'hbf, 'hbf, 'hbf, 'hbf, 'hbf, 'hbf, 'hbf,
	'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80, 'h00, 'h00, 'h00, 'h80,
	'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h00, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h81,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc7,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'hc3,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'h80, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'hc1,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'h80, 'h80, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc7, 'hc0, 'hc0, 'hc0, 'hc7, 'hc0, 'hcf, 'hcf, 'hcf,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'hc0, 'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc3,
	'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'h80, 'hc0, 'h80, 'h80, 'h80, 'hc0, 'h80, 'hc0, 'hc0, 'hc0,
	'h80, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc1,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc1, 'hc7, 'hd7,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd0, 'hc0, 'hc0, 'hc0, 'hd0, 'hc0, 'hd0, 'hd8, 'hdb,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd8,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hd8, 'hc0, 'hc0, 'hc0, 'hd8, 'hd0, 'hd8, 'hd8, 'hdd,
	'hc0, 'hc0, 'hc0, 'hd0, 'hc0, 'hd0, 'hd0, 'hdc, 'hd0, 'hd8, 'hd8, 'hdc, 'hd8, 'hdc, 'hdc, 'hde,
	'hd8, 'hdc, 'hdc, 'hde, 'hdc, 'hde, 'hde, 'hdf, 'hde, 'hdf, 'hdf, 'hdf, 'hdf, 'hdf, 'hdf, 'hdf,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he3,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'he1,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'hc0, 'hc0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'hc0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he1, 'he3, 'he7,
	'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'he0,
	'hc0, 'hc0, 'hc0, 'he0, 'hc0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'heb,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he8, 'he0, 'he8, 'he8, 'hed,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'hec, 'he0, 'he0, 'he0, 'hec, 'he8, 'hec, 'hec, 'hee,
	'he8, 'he8, 'he8, 'hec, 'hec, 'hee, 'hee, 'hef, 'hec, 'hef, 'hef, 'hef, 'hef, 'hef, 'hef, 'hef,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'hf0,
	'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'he0, 'hf0, 'he0, 'he0, 'he0, 'hf0, 'he0, 'hf0, 'hf0, 'hf0,
	'he0, 'he0, 'he0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf3,
	'he0, 'he0, 'he0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0,
	'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf5,
	'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf4, 'hf4, 'hf6,
	'hf0, 'hf0, 'hf0, 'hf4, 'hf0, 'hf4, 'hf6, 'hf7, 'hf4, 'hf6, 'hf6, 'hf7, 'hf7, 'hf7, 'hf7, 'hf7,
	'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf8, 'hf0, 'hf0, 'hf0, 'hf0, 'hf0, 'hf8, 'hf8, 'hf8,
	'hf0, 'hf0, 'hf0, 'hf8, 'hf0, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf9,
	'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hfa,
	'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hf8, 'hfb, 'hf8, 'hfa, 'hfa, 'hfb, 'hfb, 'hfb, 'hfb, 'hfb,
	'hf8, 'hf8, 'hf8, 'hfc, 'hf8, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc,
	'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfc, 'hfd, 'hfc, 'hfc, 'hfc, 'hfd, 'hfd, 'hfd, 'hfd, 'hfd,
	'hfc, 'hfc, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe, 'hfe,
	'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff, 'hff
};


/////////////////////////////////////////////////////////////////////////////////////


reg [15:0] f0;
generate
	if(MULTI_FILTERS) begin
		always_ff @(posedge ld_clk) if(ld_wr) f6581_curve[1024+ld_addr] <= ld_data;
		always_ff @(posedge clock) f0 <= f6581_curve[{cfg, Fc[10:1]}];
	end
	else begin
		always_ff @(posedge ld_clk) if(ld_wr) f6581_curve[ld_addr[9:0]] <= ld_data;
		always_ff @(posedge clock) f0 <= f6581_curve[Fc[10:1]];
	end
endgenerate

wire [10:0] fc_6581;
sid_dac #(.BITS(11)) fc_dac
(
  .vin  (Fc),
  .vout (fc_6581)
);

function reg [9:0] tanh_x_mirror(signed [10:0] x);
    tanh_x_mirror = 10'(x < 0 ? -x : x);
endfunction

function signed [10:0] tanh_x_clamp(signed [12:0] x);
    tanh_x_clamp = (x < -1023) ? -11'sd1023 :
                   (x >  1023) ?  11'sd1023 :
                   11'(x);
endfunction

function signed [15:0] tanh_y_mirror(logic x_neg,signed [15:0] y);
    tanh_y_mirror = x_neg ? -y : y;
endfunction

wire signed [15:0] f6581_adj_y0 = 16'(9883+250);
wire [10:0] fc_x = tanh_x_clamp(13'(fc_6581) - Fc_offset);

reg [15:0] f0_adj;
always_ff @(posedge clock) f0_adj <= {fc_x[10], f6581_adj[tanh_x_mirror(fc_x)]};

assign F0 = mode ? ({ 3'b000, Fc, 2'b00 } + Fc) : Fc_offset ? (f6581_adj_y0 + tanh_y_mirror(f0_adj[15], f0_adj[14:0])) : {1'b0, f0[15:1]};

// value = pi * 1.048576 * f0[fc]
reg  [15:0] f6581_curve[4*1024] =
'{
	// 0 mixed calc 
      933,    932,    932,    933,    936,    937,    943,    948,
      949,    945,    936,    926,    920,    918,    920,    924,
      930,    938,    945,    954,    960,    960,    955,    951,
      950,    949,    948,    948,    948,    945,    945,    945,
      948,    943,    942,    937,    937,    937,    939,    945,
      950,    951,    956,    960,    965,    971,    977,    981,
      982,    979,    976,    970,    964,    957,    949,    944,
      942,    942,    945,    950,    955,    955,    957,    960,
      961,    957,    954,    948,    948,    949,    955,    958,
      964,    971,    975,    979,    981,    979,    979,    975,
      973,    971,    970,    969,    969,    969,    969,    973,
      973,    971,    967,    965,    965,    963,    963,    967,
      970,    976,    987,    995,   1001,    996,    993,    987,
      983,    982,    984,    988,    992,    992,    994,    999,
      999,    994,    988,    981,    982,    988,   1002,   1014,
     1020,   1018,   1008,   1000,    994,    996,    997,   1005,
     1009,   1008,   1006,   1002,   1005,   1006,   1012,   1018,
     1024,   1024,   1024,   1024,   1026,   1027,   1029,   1033,
     1035,   1033,   1029,   1026,   1027,   1029,   1035,   1041,
     1047,   1048,   1047,   1048,   1053,   1059,   1072,   1082,
     1086,   1078,   1063,   1047,   1041,   1045,   1057,   1069,
     1078,   1082,   1086,   1087,   1090,   1090,   1089,   1087,
     1090,   1091,   1098,   1104,   1105,   1099,   1092,   1086,
     1086,   1096,   1115,   1132,   1147,   1150,   1147,   1141,
     1141,   1141,   1144,   1149,   1154,   1156,   1162,   1166,
     1174,   1180,   1187,   1194,   1197,   1193,   1189,   1183,
     1183,   1188,   1197,   1209,   1216,   1216,   1213,   1210,
     1210,   1210,   1213,   1216,   1219,   1220,   1222,   1225,
     1231,   1238,   1247,   1259,   1271,   1275,   1280,   1286,
     1293,   1297,   1303,   1306,   1310,   1308,   1306,   1306,
     1310,   1318,   1330,   1343,   1354,   1360,   1364,   1367,
     1378,   1393,   1415,   1435,   1448,   1448,   1436,   1426,
     1426,   1435,   1451,   1471,   1484,   1486,   1486,   1486,
     1490,   1498,   1510,   1520,   1535,   1545,   1555,   1564,
     1576,   1585,   1599,   1612,   1622,   1625,   1630,   1633,
     1644,   1655,   1676,   1696,   1713,   1723,   1732,   1738,
     1750,   1761,   1777,   1794,   1807,   1818,   1823,   1828,
     1840,   1857,   1880,   1904,   1921,   1931,   1937,   1944,
     1956,   1970,   1992,   2013,   2035,   2053,   2069,   2087,
     2106,   2124,   2145,   2164,   2185,   2204,   2220,   2238,
     2262,   2283,   2308,   2333,   2356,   2375,   2392,   2409,
     2429,   2448,   2468,   2488,   2510,   2537,   2567,   2601,
     2629,   2650,   2672,   2693,   2720,   2757,   2799,   2843,
     2881,   2905,   2927,   2943,   2969,   2993,   3023,   3054,
     3086,   3115,   3145,   3175,   3207,   3243,   3280,   3319,
     3353,   3385,   3415,   3444,   3472,   3493,   3511,   3531,
     3563,   3606,   3660,   3715,   3761,   3787,   3804,   3819,
     3845,   3888,   3941,   3991,   4033,   4051,   4062,   4071,
     4092,   4126,   4169,   4218,   4264,   4303,   4345,   4383,
     4424,   4460,   4493,   4530,   4575,   4629,   4692,   4755,
     4814,   4862,   4903,   4945,   4991,   5045,   5102,   5160,
     5217,   5269,   5316,   5366,   5421,   5480,   5542,   5604,
     5664,   5716,   5763,   5813,   5867,   5929,   5996,   6064,
     6129,   6185,   6240,   6294,   6354,   6415,   6483,   6548,
     6614,   6670,   6723,   6778,   6840,   6910,   6988,   7067,
     7144,   7216,   7287,   7354,   7420,   7481,   7536,   7593,
     7654,   7715,   7777,   7845,   7917,   7996,   8083,   8171,
     8255,   8332,   8408,   8482,   8558,   8628,   8696,   8768,
     8851,   8946,   9057,   9164,   9261,   9336,   9400,   9466,
     9541,   9629,   9727,   9825,   9922,  10011,  10096,  10181,
    10275,  10377,  10485,  10595,  10701,  10789,  10868,  10952,
    11056,  11187,  11336,  11485,  11617,  11719,  11803,  11886,
    11983,  12099,  12228,  12360,  12487,  12601,  12712,  12829,
    12961,  13151,  13389,  13597,  13706,  13649,  13479,  13308,
    10866,  10883,  10985,  11125,  11250,  11362,  11483,  11606,
    11720,  11813,  11899,  11984,  12076,  12180,  12294,  12408,
    12516,  12607,  12689,  12773,  12869,  12976,  13091,  13212,
    13332,  13454,  13578,  13699,  13812,  13911,  14003,  14089,
    14180,  14270,  14362,  14456,  14559,  14666,  14787,  14904,
    15011,  15096,  15172,  15250,  15344,  15458,  15590,  15723,
    15851,  15960,  16063,  16168,  16281,  16408,  16544,  16680,
    16801,  16904,  16995,  17080,  17157,  17216,  17264,  17317,
    17396,  17508,  17647,  17789,  17919,  18027,  18124,  18219,
    18315,  18410,  18504,  18601,  18705,  18821,  18944,  19070,
    19194,  19312,  19431,  19546,  19659,  19762,  19859,  19959,
    20066,  20187,  20318,  20447,  20568,  20669,  20764,  20856,
    20952,  21048,  21147,  21249,  21357,  21470,  21588,  21707,
    21828,  21951,  22076,  22197,  22316,  22424,  22528,  22631,
    22743,  22864,  22992,  23120,  23247,  23367,  23484,  23602,
    23725,  23869,  24031,  24170,  24251,  24230,  24142,  24052,
    24037,  24125,  24274,  24443,  24594,  24714,  24827,  24937,
    25049,  25168,  25289,  25406,  25517,  25609,  25693,  25777,
    25879,  26004,  26147,  26290,  26416,  26514,  26599,  26682,
    26781,  26908,  27050,  27190,  27308,  27392,  27454,  27517,
    27599,  27712,  27845,  27978,  28094,  28181,  28248,  28319,
    28412,  28541,  28691,  28841,  28968,  29059,  29133,  29201,
    29281,  29375,  29476,  29582,  29688,  29797,  29910,  30022,
    30130,  30229,  30326,  30419,  30505,  30578,  30643,  30707,
    30781,  30867,  30960,  31056,  31146,  31228,  31308,  31386,
    31467,  31551,  31635,  31722,  31813,  31904,  31998,  32093,
    32192,  32292,  32395,  32496,  32591,  32674,  32750,  32825,
    32911,  33009,  33116,  33222,  33313,  33383,  33440,  33497,
    33566,  33654,  33752,  33851,  33941,  34014,  34078,  34139,
    34205,  34273,  34344,  34415,  34487,  34559,  34632,  34705,
    34773,  34832,  34888,  34942,  35004,  35073,  35146,  35220,
    35292,  35371,  35458,  35526,  35552,  35506,  35408,  35310,
    35265,  35298,  35375,  35468,  35544,  35594,  35636,  35677,
    35727,  35788,  35855,  35922,  35982,  36033,  36079,  36121,
    36159,  36187,  36207,  36231,  36269,  36327,  36399,  36473,
    36540,  36601,  36659,  36710,  36751,  36771,  36778,  36785,
    36806,  36846,  36899,  36954,  37004,  37047,  37088,  37125,
    37157,  37182,  37200,  37218,  37243,  37276,  37312,  37352,
    37390,  37427,  37466,  37504,  37540,  37574,  37607,  37640,
    37672,  37708,  37745,  37780,  37809,  37829,  37843,  37857,
    37874,  37893,  37914,  37937,  37962,  37992,  38024,  38057,
    38090,  38120,  38151,  38181,  38210,  38238,  38267,  38294,
    38318,  38340,  38359,  38378,  38398,  38418,  38438,  38459,
    38480,  38502,  38525,  38548,  38569,  38590,  38609,  38627,
    38646,  38665,  38685,  38704,  38723,  38742,  38761,  38780,
    38798,  38817,  38837,  38855,  38870,  38880,  38887,  38895,
    38905,  38920,  38937,  38954,  38973,  38992,  39013,  39032,
    39047,  39058,  39065,  39070,  39072,  39071,  39066,  39061,
    39061,  39064,  39070,  39079,  39088,  39099,  39112,  39125,
    39136,  39142,  39143,  39145,  39146,  39148,  39149,  39151,
    39152,  39154,  39155,  39156,  39158,  39159,  39160,  39161,
    39163,  39164,  39165,  39166,  39168,  39169,  39170,  39171,
    39172,  39173,  39174,  39175,  39176,  39177,  39178,  39179,
    39180,  39181,  39182,  39183,  39184,  39185,  39186,  39187,
    39188,  39189,  39189,  39190,  39191,  39192,  39193,  39194,
    39194,  39195,  39196,  39197,  39198,  39198,  39199,  39200,
    39201,  39202,  39202,  39203,  39204,  39204,  39205,  39206,
    39207,  39207,  39208,  39209,  39209,  39210,  39210,  39211,
    39212,  39212,  39213,  39213,  39214,  39214,  39215,  39215,
    39216,  39216,  39217,  39217,  39218,  39218,  39219,  39219,
    39220,  39220,  39220,  39221,  39221,  39222,  39222,  39222,
    39223,  39223,  39224,  39224,  39224,  39225,  39225,  39226,
    39226,  39226,  39227,  39227,  39227,  39228,  39228,  39228,
    39229,  39229,  39229,  39230,  39230,  39231,  39231,  39231,
	 

	// 1 web 
      843,    840,    840,    843,    846,    849,    859,    866,
      869,    859,    843,    826,    816,    813,    816,    823,
      833,    843,    856,    869,    879,    879,    872,    866,
      863,    859,    856,    856,    856,    853,    853,    853,
      853,    846,    843,    836,    836,    836,    840,    846,
      853,    856,    863,    869,    879,    886,    896,    902,
      905,    899,    892,    882,    872,    859,    846,    833,
      830,    830,    836,    843,    849,    849,    853,    856,
      856,    849,    843,    833,    833,    833,    843,    849,
      859,    866,    872,    879,    882,    879,    876,    869,
      866,    863,    859,    856,    856,    856,    856,    859,
      859,    856,    849,    843,    843,    840,    840,    843,
      849,    859,    872,    886,    896,    889,    879,    869,
      863,    859,    863,    869,    872,    872,    876,    879,
      879,    869,    859,    846,    846,    856,    876,    896,
      905,    899,    882,    866,    856,    856,    859,    866,
      872,    869,    863,    856,    856,    859,    866,    876,
      882,    882,    879,    879,    879,    879,    882,    886,
      889,    882,    876,    866,    866,    869,    876,    886,
      892,    892,    889,    889,    892,    902,    922,    935,
      942,    925,    896,    869,    856,    859,    876,    896,
      909,    912,    915,    915,    915,    912,    909,    905,
      905,    905,    912,    919,    919,    905,    889,    872,
      869,    882,    912,    938,    958,    958,    948,    935,
      928,    925,    928,    932,    935,    935,    942,    945,
      952,    958,    968,    975,    978,    968,    955,    942,
      938,    942,    955,    968,    978,    975,    965,    955,
      952,    948,    948,    948,    948,    945,    945,    942,
      948,    955,    968,    981,    994,    998,   1001,   1004,
     1008,   1008,   1011,   1011,   1011,   1001,    991,    981,
      981,    988,    998,   1014,   1024,   1024,   1021,   1017,
     1024,   1040,   1067,   1090,   1103,   1090,   1060,   1031,
     1017,   1021,   1037,   1057,   1067,   1060,   1047,   1034,
     1027,   1027,   1034,   1040,   1050,   1054,   1057,   1060,
     1067,   1070,   1080,   1087,   1090,   1083,   1073,   1067,
     1067,   1073,   1093,   1110,   1123,   1123,   1123,   1116,
     1120,   1123,   1133,   1143,   1149,   1146,   1136,   1129,
     1129,   1139,   1156,   1176,   1185,   1182,   1169,   1159,
     1156,   1159,   1172,   1185,   1199,   1202,   1208,   1212,
     1218,   1222,   1232,   1238,   1245,   1248,   1248,   1251,
     1258,   1264,   1278,   1288,   1297,   1297,   1294,   1291,
     1291,   1288,   1288,   1288,   1294,   1304,   1320,   1340,
     1353,   1353,   1350,   1350,   1360,   1383,   1419,   1456,
     1482,   1485,   1479,   1469,   1469,   1472,   1482,   1492,
     1505,   1512,   1521,   1531,   1544,   1561,   1581,   1604,
     1620,   1630,   1637,   1640,   1643,   1633,   1617,   1604,
     1610,   1640,   1686,   1736,   1765,   1762,   1742,   1719,
     1716,   1739,   1782,   1821,   1841,   1824,   1792,   1755,
     1739,   1745,   1768,   1798,   1821,   1831,   1841,   1848,
     1854,   1851,   1844,   1841,   1851,   1877,   1917,   1956,
     1986,   1996,   1992,   1992,   1999,   2016,   2039,   2062,
     2085,   2095,   2101,   2108,   2124,   2147,   2177,   2207,
     2233,   2243,   2246,   2253,   2266,   2292,   2328,   2365,
     2394,   2411,   2421,   2431,   2447,   2470,   2500,   2529,
     2556,   2566,   2569,   2576,   2595,   2628,   2674,   2724,
     2767,   2800,   2833,   2859,   2882,   2892,   2895,   2898,
     2908,   2918,   2931,   2951,   2981,   3024,   3076,   3136,
     3185,   3221,   3254,   3287,   3317,   3340,   3356,   3379,
     3422,   3491,   3584,   3673,   3742,   3771,   3778,   3785,
     3811,   3860,   3929,   3999,   4065,   4114,   4157,   4200,
     4256,   4328,   4410,   4493,   4562,   4595,   4608,   4628,
     4684,   4793,   4938,   5082,   5194,   5244,   5260,   5270,
     5313,   5395,   5501,   5610,   5708,   5774,   5827,   5886,
     5969,   6143,   6384,   6548,   6506,   6117,   5488,   4849,
     4420,   4282,   4312,   4420,   4516,   4595,   4697,   4802,
     4891,   4941,   4977,   5010,   5059,   5135,   5227,   5320,
     5395,   5438,   5461,   5488,   5534,   5606,   5692,   5791,
     5890,   5992,   6100,   6206,   6295,   6357,   6407,   6450,
     6502,   6558,   6621,   6690,   6776,   6881,   7010,   7135,
     7240,   7303,   7342,   7388,   7467,   7593,   7754,   7919,
     8067,   8182,   8281,   8383,   8505,   8657,   8831,   9003,
     9144,   9246,   9325,   9388,   9437,   9447,   9431,   9427,
     9480,   9615,   9806,  10007,  10182,  10307,  10409,  10505,
    10607,  10706,  10804,  10907,  11032,  11180,  11348,  11523,
    11694,  11852,  12013,  12168,  12317,  12442,  12557,  12676,
    12814,  12985,  13183,  13377,  13549,  13680,  13792,  13898,
    14013,  14135,  14260,  14392,  14540,  14702,  14876,  15057,
    15242,  15430,  15624,  15815,  15996,  16154,  16299,  16444,
    16612,  16803,  17014,  17228,  17439,  17630,  17818,  18006,
    18210,  18473,  18783,  19033,  19129,  18951,  18589,  18226,
    18062,  18174,  18450,  18786,  19070,  19271,  19455,  19633,
    19817,  20018,  20229,  20433,  20615,  20750,  20858,  20970,
    21132,  21362,  21646,  21929,  22166,  22324,  22443,  22558,
    22723,  22967,  23260,  23550,  23777,  23899,  23958,  24018,
    24139,  24357,  24634,  24917,  25147,  25286,  25368,  25460,
    25625,  25902,  26251,  26603,  26883,  27051,  27160,  27256,
    27387,  27569,  27773,  27997,  28224,  28461,  28715,  28969,
    29206,  29423,  29631,  29825,  29996,  30125,  30227,  30326,
    30461,  30639,  30846,  31064,  31261,  31429,  31588,  31746,
    31914,  32092,  32276,  32470,  32678,  32892,  33119,  33353,
    33597,  33854,  34124,  34391,  34635,  34832,  35004,  35178,
    35389,  35659,  35972,  36279,  36532,  36694,  36802,  36911,
    37076,  37326,  37626,  37935,  38199,  38397,  38558,  38706,
    38878,  39065,  39266,  39471,  39681,  39899,  40126,  40350,
    40558,  40729,  40881,  41032,  41220,  41447,  41704,  41968,
    42225,  42528,  42870,  43124,  43154,  42798,  42172,  41553,
    41213,  41279,  41589,  41977,  42284,  42458,  42590,  42719,
    42897,  43140,  43427,  43714,  43967,  44171,  44349,  44507,
    44642,  44722,  44758,  44817,  44962,  45229,  45585,  45960,
    46299,  46603,  46899,  47153,  47340,  47400,  47370,  47340,
    47403,  47597,  47877,  48177,  48444,  48668,  48882,  49073,
    49235,  49340,  49403,  49465,  49574,  49742,  49946,  50167,
    50388,  50605,  50829,  51056,  51274,  51475,  51669,  51863,
    52064,  52288,  52529,  52753,  52931,  53036,  53095,  53145,
    53221,  53323,  53441,  53576,  53741,  53939,  54169,  54410,
    54647,  54874,  55102,  55329,  55553,  55774,  55998,  56212,
    56406,  56571,  56712,  56851,  57002,  57160,  57322,  57493,
    57674,  57869,  58076,  58287,  58488,  58672,  58847,  59022,
    59206,  59394,  59588,  59786,  59987,  60188,  60395,  60606,
    60817,  61041,  61275,  61496,  61677,  61785,  61848,  61914,
    62033,  62217,  62448,  62701,  62971,  63274,  63614,  63933,
    64180,  64342,  64447,  64500,  64510,  64434,  64292,  64147,
    64085,  64114,  64200,  64329,  64490,  64694,  64948,  65208,
    65439,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
    65535,  65535,  65535,  65535,  65535,  65535,  65535,  65535,
	 
	 
	 
	// 2 resid 6581
      724,    724,    724,    724,    724,    724,    724,    724,
      724,    728,    728,    728,    728,    728,    728,    728,
      728,    731,    731,    731,    731,    731,    731,    731,
      731,    734,    734,    734,    734,    734,    734,    734,
      737,    737,    737,    737,    737,    737,    737,    741,
      741,    741,    741,    741,    741,    744,    744,    744,
      744,    744,    747,    747,    747,    747,    747,    751,
      751,    751,    751,    751,    754,    754,    754,    754,
      757,    757,    757,    757,    757,    760,    760,    760,
      760,    764,    764,    764,    764,    764,    767,    767,
      767,    767,    770,    770,    770,    770,    770,    774,
      774,    774,    774,    777,    777,    777,    777,    780,
      780,    780,    784,    784,    784,    784,    787,    787,
      787,    790,    790,    790,    793,    793,    793,    797,
      797,    800,    800,    800,    803,    803,    807,    807,
      807,    810,    810,    813,    813,    816,    816,    820,
      823,    823,    826,    826,    830,    830,    833,    833,
      836,    836,    840,    840,    843,    846,    846,    849,
      849,    853,    853,    856,    859,    859,    863,    863,
      866,    869,    869,    872,    876,    876,    879,    882,
      882,    886,    889,    889,    892,    896,    899,    899,
      902,    905,    909,    912,    915,    919,    919,    922,
      925,    928,    932,    935,    938,    942,    945,    952,
      955,    958,    961,    965,    968,    975,    978,    981,
      988,    991,    994,    998,   1004,   1008,   1011,   1014,
     1021,   1024,   1027,   1031,   1034,   1037,   1044,   1047,
     1050,   1054,   1057,   1064,   1067,   1070,   1073,   1080,
     1083,   1087,   1090,   1096,   1100,   1106,   1110,   1116,
     1120,   1126,   1129,   1136,   1143,   1146,   1152,   1159,
     1166,   1172,   1179,   1185,   1192,   1199,   1205,   1215,
     1222,   1228,   1238,   1245,   1255,   1264,   1274,   1284,
     1294,   1304,   1314,   1324,   1334,   1347,   1357,   1370,
     1383,   1393,   1406,   1419,   1432,   1442,   1456,   1469,
     1482,   1495,   1508,   1521,   1535,   1548,   1561,   1574,
     1587,   1600,   1614,   1630,   1643,   1656,   1673,   1686,
     1703,   1716,   1732,   1749,   1765,   1782,   1798,   1815,
     1831,   1848,   1864,   1884,   1900,   1920,   1940,   1956,
     1976,   1996,   2016,   2039,   2058,   2078,   2101,   2124,
     2147,   2167,   2193,   2216,   2240,   2266,   2289,   2315,
     2342,   2368,   2394,   2421,   2450,   2480,   2506,   2536,
     2569,   2599,   2628,   2661,   2691,   2724,   2757,   2790,
     2823,   2859,   2892,   2928,   2961,   2997,   3033,   3070,
     3106,   3142,   3182,   3218,   3257,   3297,   3333,   3373,
     3412,   3452,   3495,   3534,   3577,   3617,   3659,   3702,
     3745,   3788,   3831,   3873,   3916,   3962,   4005,   4051,
     4094,   4140,   4186,   4233,   4279,   4325,   4374,   4420,
     4470,   4516,   4565,   4611,   4661,   4710,   4760,   4809,
     4858,   4911,   4961,   5010,   5063,   5112,   5165,   5218,
     5270,   5323,   5376,   5432,   5491,   5550,   5613,   5675,
     5741,   5807,   5873,   5942,   6011,   6081,   6153,   6226,
     6301,   6377,   6453,   6529,   6604,   6683,   6762,   6842,
     6921,   7003,   7082,   7164,   7247,   7329,   7411,   7494,
     7576,   7659,   7741,   7823,   7909,   7995,   8080,   8166,
     8255,   8340,   8429,   8518,   8611,   8699,   8792,   8881,
     8976,   9068,   9161,   9256,   9352,   9447,   9543,   9638,
     9737,   9836,   9935,  10034,  10132,  10235,  10333,  10436,
    10541,  10643,  10745,  10851,  10956,  11061,  11170,  11276,
    11384,  11493,  11602,  11710,  11822,  11931,  12043,  12155,
    12270,  12382,  12498,  12613,  12728,  12844,  12959,  13077,
    13196,  13315,  13433,  13552,  13674,  13796,  13917,  14039,
    14165,  14290,  14418,  14550,  14688,  14827,  14968,  15113,
    15262,  15410,  15558,  15710,  15861,  16013,  16164,  16319,
    16470,  16619,  16774,  16928,  17087,  17251,  17423,  17600,
    17788,  17999,  18246,  18510,  18776,  19047,  19327,  19616,
    15153,  15324,  15495,  15660,  15812,  15953,  16092,  16230,
    16368,  16503,  16638,  16774,  16909,  17044,  17179,  17317,
    17459,  17600,  17742,  17887,  18035,  18180,  18328,  18477,
    18625,  18773,  18918,  19063,  19208,  19350,  19491,  19626,
    19765,  19896,  20025,  20153,  20282,  20404,  20529,  20651,
    20773,  20891,  21013,  21132,  21254,  21372,  21494,  21616,
    21741,  21863,  21988,  22113,  22235,  22361,  22486,  22611,
    22736,  22861,  22983,  23108,  23230,  23352,  23474,  23596,
    23718,  23836,  23955,  24074,  24192,  24311,  24429,  24548,
    24666,  24782,  24900,  25019,  25134,  25253,  25371,  25487,
    25605,  25721,  25839,  25954,  26070,  26188,  26304,  26422,
    26538,  26656,  26771,  26887,  27005,  27121,  27239,  27355,
    27473,  27588,  27704,  27822,  27941,  28056,  28175,  28290,
    28409,  28527,  28646,  28761,  28880,  28998,  29117,  29236,
    29354,  29476,  29595,  29713,  29832,  29954,  30072,  30194,
    30316,  30435,  30556,  30678,  30800,  30922,  31047,  31169,
    31294,  31416,  31541,  31663,  31789,  31914,  32039,  32164,
    32289,  32418,  32543,  32668,  32797,  32922,  33050,  33179,
    33304,  33432,  33561,  33689,  33818,  33946,  34075,  34203,
    34332,  34463,  34592,  34720,  34849,  34981,  35109,  35241,
    35369,  35498,  35630,  35758,  35890,  36022,  36150,  36282,
    36410,  36542,  36671,  36802,  36934,  37063,  37194,  37323,
    37455,  37583,  37715,  37843,  37975,  38103,  38235,  38364,
    38496,  38624,  38752,  38884,  39013,  39141,  39270,  39398,
    39530,  39658,  39787,  39919,  40050,  40182,  40314,  40446,
    40581,  40716,  40848,  40983,  41121,  41256,  41391,  41526,
    41665,  41800,  41938,  42076,  42211,  42350,  42488,  42623,
    42761,  42900,  43035,  43173,  43308,  43443,  43582,  43717,
    43852,  43987,  44122,  44254,  44389,  44521,  44652,  44784,
    44916,  45048,  45176,  45305,  45433,  45562,  45687,  45812,
    45937,  46059,  46181,  46303,  46425,  46543,  46659,  46777,
    46892,  47004,  47120,  47228,  47340,  47449,  47555,  47660,
    47765,  47868,  47966,  48068,  48164,  48263,  48358,  48454,
    48549,  48642,  48734,  48823,  48912,  49001,  49090,  49175,
    49261,  49347,  49429,  49515,  49597,  49676,  49758,  49837,
    49916,  49996,  50071,  50147,  50223,  50299,  50374,  50450,
    50523,  50595,  50668,  50740,  50813,  50882,  50954,  51023,
    51093,  51162,  51231,  51300,  51369,  51438,  51504,  51573,
    51639,  51705,  51774,  51840,  51906,  51972,  52041,  52107,
    52173,  52239,  52305,  52371,  52440,  52506,  52572,  52638,
    52707,  52773,  52838,  52904,  52970,  53036,  53102,  53168,
    53234,  53296,  53362,  53425,  53491,  53553,  53616,  53678,
    53741,  53804,  53866,  53929,  53991,  54051,  54113,  54173,
    54232,  54291,  54354,  54410,  54469,  54528,  54588,  54644,
    54703,  54759,  54815,  54871,  54927,  54983,  55039,  55095,
    55148,  55204,  55256,  55309,  55362,  55415,  55467,  55517,
    55569,  55619,  55671,  55721,  55770,  55820,  55869,  55915,
    55965,  56011,  56057,  56103,  56149,  56195,  56241,  56284,
    56330,  56373,  56416,  56459,  56498,  56541,  56581,  56620,
    56660,  56699,  56739,  56778,  56815,  56851,  56890,  56927,
    56963,  56996,  57032,  57068,  57101,  57134,  57167,  57200,
    57233,  57266,  57299,  57328,  57361,  57391,  57421,  57450,
    57480,  57510,  57539,  57569,  57595,  57625,  57651,  57681,
    57707,  57734,  57763,  57790,  57816,  57842,  57869,  57892,
    57918,  57944,  57968,  57994,  58017,  58043,  58066,  58093,
    58116,  58139,  58165,  58188,  58211,  58234,  58257,  58280,
    58307,  58330,  58350,  58373,  58396,  58416,  58439,  58458,
    58481,  58501,  58521,  58541,  58560,  58580,  58597,  58616,
    58636,  58653,  58669,  58689,  58705,  58722,  58738,  58755,
    58771,  58788,  58804,  58821,  58834,  58850,  58864,  58880,
    58893,  58910,  58923,  58936,  58952,  58966,  58979,  58992,
    59005,  59018,  59032,  59045,  59058,  59071,  59084,  59097,
    59107,  59120,  59134,  59144,  59157,  59170,  59180,  59193,
    59206,  59216,  59229,  59239,  59252,  59265,  59275,  59288,
	 
	 

	// 3 resid 6581/2
      362,    362,    362,    362,    362,    362,    362,    362,
      362,    364,    364,    364,    364,    364,    364,    364,
      364,    365,    365,    365,    365,    365,    365,    365,
      365,    367,    367,    367,    367,    367,    367,    367,
      368,    368,    368,    368,    368,    368,    368,    370,
      370,    370,    370,    370,    370,    372,    372,    372,
      372,    372,    373,    373,    373,    373,    373,    375,
      375,    375,    375,    375,    377,    377,    377,    377,
      378,    378,    378,    378,    378,    380,    380,    380,
      380,    382,    382,    382,    382,    382,    383,    383,
      383,    383,    385,    385,    385,    385,    385,    387,
      387,    387,    387,    388,    388,    388,    388,    390,
      390,    390,    392,    392,    392,    392,    393,    393,
      393,    395,    395,    395,    396,    396,    396,    398,
      398,    400,    400,    400,    401,    401,    403,    403,
      403,    405,    405,    406,    406,    408,    408,    410,
      411,    411,    413,    413,    415,    415,    416,    416,
      418,    418,    420,    420,    421,    423,    423,    424,
      424,    426,    426,    428,    429,    429,    431,    431,
      433,    434,    434,    436,    438,    438,    439,    441,
      441,    443,    444,    444,    446,    448,    449,    449,
      451,    452,    454,    456,    457,    459,    459,    461,
      462,    464,    466,    467,    469,    471,    472,    476,
      477,    479,    480,    482,    484,    487,    489,    490,
      494,    495,    497,    499,    502,    504,    505,    507,
      510,    512,    513,    515,    517,    518,    522,    523,
      525,    527,    528,    532,    533,    535,    536,    540,
      541,    543,    545,    548,    550,    553,    555,    558,
      560,    563,    564,    568,    571,    573,    576,    579,
      583,    586,    589,    592,    596,    599,    602,    607,
      611,    614,    619,    622,    627,    632,    637,    642,
      647,    652,    657,    662,    667,    673,    678,    685,
      691,    696,    703,    709,    716,    721,    728,    734,
      741,    747,    754,    760,    767,    774,    780,    787,
      793,    800,    807,    815,    821,    828,    836,    843,
      851,    858,    866,    874,    882,    891,    899,    907,
      915,    924,    932,    942,    950,    960,    970,    978,
      988,    998,   1008,   1019,   1029,   1039,   1050,   1062,
     1073,   1083,   1096,   1108,   1120,   1133,   1144,   1157,
     1171,   1184,   1197,   1210,   1225,   1240,   1253,   1268,
     1284,   1299,   1314,   1330,   1345,   1362,   1378,   1395,
     1411,   1429,   1446,   1464,   1480,   1498,   1516,   1535,
     1553,   1571,   1591,   1609,   1628,   1648,   1666,   1686,
     1706,   1726,   1747,   1767,   1788,   1808,   1829,   1851,
     1872,   1894,   1915,   1936,   1958,   1981,   2002,   2025,
     2047,   2070,   2093,   2116,   2139,   2162,   2187,   2210,
     2235,   2258,   2282,   2305,   2330,   2355,   2380,   2404,
     2429,   2455,   2480,   2505,   2531,   2556,   2582,   2609,
     2635,   2661,   2688,   2716,   2745,   2775,   2806,   2837,
     2870,   2903,   2936,   2971,   3005,   3040,   3076,   3113,
     3150,   3188,   3226,   3264,   3302,   3341,   3381,   3421,
     3460,   3501,   3541,   3582,   3623,   3664,   3705,   3747,
     3788,   3829,   3870,   3911,   3954,   3997,   4040,   4083,
     4127,   4170,   4214,   4259,   4305,   4349,   4396,   4440,
     4488,   4534,   4580,   4628,   4676,   4723,   4771,   4819,
     4868,   4918,   4967,   5017,   5066,   5117,   5166,   5218,
     5270,   5321,   5372,   5425,   5478,   5530,   5585,   5638,
     5692,   5746,   5801,   5855,   5911,   5965,   6021,   6077,
     6135,   6191,   6249,   6306,   6364,   6422,   6479,   6538,
     6598,   6657,   6716,   6776,   6837,   6898,   6958,   7019,
     7082,   7145,   7209,   7275,   7344,   7413,   7484,   7556,
     7631,   7705,   7779,   7855,   7930,   8006,   8082,   8159,
     8235,   8309,   8387,   8464,   8543,   8625,   8711,   8800,
     8894,   8999,   9123,   9255,   9388,   9523,   9663,   9808,
     7576,   7662,   7747,   7830,   7906,   7976,   8046,   8115,
     8184,   8251,   8319,   8387,   8454,   8522,   8589,   8658,
     8729,   8800,   8871,   8943,   9017,   9090,   9164,   9238,
     9312,   9386,   9459,   9531,   9604,   9675,   9745,   9813,
     9882,   9948,  10012,  10076,  10141,  10202,  10264,  10325,
    10386,  10445,  10506,  10566,  10627,  10686,  10747,  10808,
    10870,  10931,  10994,  11056,  11117,  11180,  11243,  11305,
    11368,  11430,  11491,  11554,  11615,  11676,  11737,  11798,
    11859,  11918,  11977,  12037,  12096,  12155,  12214,  12274,
    12333,  12391,  12450,  12509,  12567,  12626,  12685,  12743,
    12802,  12860,  12919,  12977,  13035,  13094,  13152,  13211,
    13269,  13328,  13385,  13443,  13502,  13560,  13619,  13677,
    13736,  13794,  13852,  13911,  13970,  14028,  14087,  14145,
    14204,  14263,  14323,  14380,  14440,  14499,  14558,  14618,
    14677,  14738,  14797,  14856,  14916,  14977,  15036,  15097,
    15158,  15217,  15278,  15339,  15400,  15461,  15523,  15584,
    15647,  15708,  15770,  15831,  15894,  15957,  16019,  16082,
    16144,  16209,  16271,  16334,  16398,  16461,  16525,  16589,
    16652,  16716,  16780,  16844,  16909,  16973,  17037,  17101,
    17166,  17231,  17296,  17360,  17424,  17490,  17554,  17620,
    17684,  17749,  17815,  17879,  17945,  18011,  18075,  18141,
    18205,  18271,  18335,  18401,  18467,  18531,  18597,  18661,
    18727,  18791,  18857,  18921,  18987,  19051,  19117,  19182,
    19248,  19312,  19376,  19442,  19506,  19570,  19635,  19699,
    19765,  19829,  19893,  19959,  20025,  20091,  20157,  20223,
    20290,  20358,  20424,  20491,  20560,  20628,  20695,  20763,
    20832,  20900,  20969,  21038,  21105,  21175,  21244,  21311,
    21380,  21450,  21517,  21586,  21654,  21721,  21791,  21858,
    21926,  21993,  22061,  22127,  22194,  22260,  22326,  22392,
    22458,  22524,  22588,  22652,  22716,  22781,  22843,  22906,
    22968,  23029,  23090,  23151,  23212,  23271,  23329,  23388,
    23446,  23502,  23560,  23614,  23670,  23724,  23777,  23830,
    23882,  23934,  23983,  24034,  24082,  24131,  24179,  24227,
    24274,  24321,  24367,  24411,  24456,  24500,  24545,  24587,
    24630,  24673,  24714,  24757,  24798,  24838,  24879,  24918,
    24958,  24998,  25035,  25073,  25111,  25149,  25187,  25225,
    25261,  25297,  25334,  25370,  25406,  25441,  25477,  25511,
    25546,  25581,  25615,  25650,  25684,  25719,  25752,  25786,
    25819,  25852,  25887,  25920,  25953,  25986,  26020,  26053,
    26086,  26119,  26152,  26185,  26220,  26253,  26286,  26319,
    26353,  26386,  26419,  26452,  26485,  26518,  26551,  26584,
    26617,  26648,  26681,  26712,  26745,  26776,  26808,  26839,
    26870,  26902,  26933,  26964,  26995,  27025,  27056,  27086,
    27116,  27145,  27177,  27205,  27234,  27264,  27294,  27322,
    27351,  27379,  27407,  27435,  27463,  27491,  27519,  27547,
    27574,  27602,  27628,  27654,  27681,  27707,  27733,  27758,
    27784,  27809,  27835,  27860,  27885,  27910,  27934,  27957,
    27982,  28005,  28028,  28051,  28074,  28097,  28120,  28142,
    28165,  28186,  28208,  28229,  28249,  28270,  28290,  28310,
    28330,  28349,  28369,  28389,  28407,  28425,  28445,  28463,
    28481,  28498,  28516,  28534,  28550,  28567,  28583,  28600,
    28616,  28633,  28649,  28664,  28680,  28695,  28710,  28725,
    28740,  28755,  28769,  28784,  28797,  28812,  28825,  28840,
    28853,  28867,  28881,  28895,  28908,  28921,  28934,  28946,
    28959,  28972,  28984,  28997,  29008,  29021,  29033,  29046,
    29058,  29069,  29082,  29094,  29105,  29117,  29128,  29140,
    29153,  29165,  29175,  29186,  29198,  29208,  29219,  29229,
    29240,  29250,  29260,  29270,  29280,  29290,  29298,  29308,
    29318,  29326,  29334,  29344,  29352,  29361,  29369,  29377,
    29385,  29394,  29402,  29410,  29417,  29425,  29432,  29440,
    29446,  29455,  29461,  29468,  29476,  29483,  29489,  29496,
    29502,  29509,  29516,  29522,  29529,  29535,  29542,  29548,
    29553,  29560,  29567,  29572,  29578,  29585,  29590,  29596,
    29603,  29608,  29614,  29619,  29626,  29632,  29637,  29644
};

//reDIP-SID curve
wire [14:0] f6581_adj[1024] =
'{
       0,     28,     56,     85,    113,    141,    169,    198,
     226,    254,    282,    310,    339,    367,    395,    423,
     451,    480,    508,    536,    564,    592,    620,    648,
     677,    705,    733,    761,    789,    817,    845,    873,
     901,    929,    957,    985,   1013,   1041,   1069,   1097,
    1125,   1152,   1180,   1208,   1236,   1264,   1291,   1319,
    1347,   1375,   1402,   1430,   1458,   1485,   1513,   1540,
    1568,   1595,   1623,   1650,   1678,   1705,   1733,   1760,
    1787,   1815,   1842,   1869,   1896,   1923,   1951,   1978,
    2005,   2032,   2059,   2086,   2113,   2140,   2167,   2194,
    2220,   2247,   2274,   2301,   2327,   2354,   2381,   2407,
    2434,   2460,   2487,   2513,   2539,   2566,   2592,   2618,
    2645,   2671,   2697,   2723,   2749,   2775,   2801,   2827,
    2853,   2879,   2905,   2931,   2956,   2982,   3008,   3033,
    3059,   3084,   3110,   3135,   3160,   3186,   3211,   3236,
    3262,   3287,   3312,   3337,   3362,   3387,   3412,   3436,
    3461,   3486,   3511,   3535,   3560,   3584,   3609,   3633,
    3658,   3682,   3706,   3731,   3755,   3779,   3803,   3827,
    3851,   3875,   3899,   3923,   3946,   3970,   3994,   4017,
    4041,   4064,   4088,   4111,   4135,   4158,   4181,   4204,
    4227,   4250,   4273,   4296,   4319,   4342,   4365,   4387,
    4410,   4433,   4455,   4478,   4500,   4522,   4545,   4567,
    4589,   4611,   4633,   4655,   4677,   4699,   4721,   4743,
    4764,   4786,   4808,   4829,   4851,   4872,   4893,   4915,
    4936,   4957,   4978,   4999,   5020,   5041,   5062,   5083,
    5103,   5124,   5145,   5165,   5186,   5206,   5227,   5247,
    5267,   5287,   5307,   5328,   5348,   5367,   5387,   5407,
    5427,   5447,   5466,   5486,   5505,   5525,   5544,   5563,
    5583,   5602,   5621,   5640,   5659,   5678,   5697,   5716,
    5734,   5753,   5772,   5790,   5809,   5827,   5846,   5864,
    5882,   5901,   5919,   5937,   5955,   5973,   5991,   6008,
    6026,   6044,   6062,   6079,   6097,   6114,   6132,   6149,
    6166,   6183,   6200,   6218,   6235,   6252,   6268,   6285,
    6302,   6319,   6336,   6352,   6369,   6385,   6402,   6418,
    6434,   6450,   6467,   6483,   6499,   6515,   6531,   6547,
    6562,   6578,   6594,   6609,   6625,   6641,   6656,   6671,
    6687,   6702,   6717,   6732,   6748,   6763,   6778,   6793,
    6807,   6822,   6837,   6852,   6866,   6881,   6895,   6910,
    6924,   6939,   6953,   6967,   6981,   6995,   7009,   7023,
    7037,   7051,   7065,   7079,   7093,   7106,   7120,   7133,
    7147,   7160,   7174,   7187,   7200,   7214,   7227,   7240,
    7253,   7266,   7279,   7292,   7305,   7317,   7330,   7343,
    7355,   7368,   7380,   7393,   7405,   7418,   7430,   7442,
    7454,   7467,   7479,   7491,   7503,   7515,   7527,   7538,
    7550,   7562,   7574,   7585,   7597,   7608,   7620,   7631,
    7643,   7654,   7665,   7676,   7688,   7699,   7710,   7721,
    7732,   7743,   7754,   7764,   7775,   7786,   7797,   7807,
    7818,   7828,   7839,   7849,   7860,   7870,   7880,   7891,
    7901,   7911,   7921,   7931,   7941,   7951,   7961,   7971,
    7981,   7991,   8000,   8010,   8020,   8029,   8039,   8049,
    8058,   8067,   8077,   8086,   8096,   8105,   8114,   8123,
    8132,   8141,   8150,   8159,   8168,   8177,   8186,   8195,
    8204,   8213,   8221,   8230,   8239,   8247,   8256,   8264,
    8273,   8281,   8290,   8298,   8306,   8315,   8323,   8331,
    8339,   8347,   8355,   8363,   8371,   8379,   8387,   8395,
    8403,   8411,   8418,   8426,   8434,   8442,   8449,   8457,
    8464,   8472,   8479,   8487,   8494,   8501,   8509,   8516,
    8523,   8531,   8538,   8545,   8552,   8559,   8566,   8573,
    8580,   8587,   8594,   8601,   8608,   8614,   8621,   8628,
    8635,   8641,   8648,   8654,   8661,   8668,   8674,   8681,
    8687,   8693,   8700,   8706,   8712,   8719,   8725,   8731,
    8737,   8743,   8750,   8756,   8762,   8768,   8774,   8780,
    8786,   8792,   8797,   8803,   8809,   8815,   8821,   8826,
    8832,   8838,   8843,   8849,   8855,   8860,   8866,   8871,
    8877,   8882,   8887,   8893,   8898,   8904,   8909,   8914,
    8919,   8925,   8930,   8935,   8940,   8945,   8950,   8955,
    8960,   8965,   8970,   8975,   8980,   8985,   8990,   8995,
    9000,   9005,   9009,   9014,   9019,   9024,   9028,   9033,
    9038,   9042,   9047,   9051,   9056,   9060,   9065,   9069,
    9074,   9078,   9083,   9087,   9091,   9096,   9100,   9104,
    9108,   9113,   9117,   9121,   9125,   9129,   9134,   9138,
    9142,   9146,   9150,   9154,   9158,   9162,   9166,   9170,
    9174,   9178,   9181,   9185,   9189,   9193,   9197,   9201,
    9204,   9208,   9212,   9215,   9219,   9223,   9226,   9230,
    9234,   9237,   9241,   9244,   9248,   9251,   9255,   9258,
    9262,   9265,   9269,   9272,   9275,   9279,   9282,   9285,
    9289,   9292,   9295,   9298,   9302,   9305,   9308,   9311,
    9314,   9318,   9321,   9324,   9327,   9330,   9333,   9336,
    9339,   9342,   9345,   9348,   9351,   9354,   9357,   9360,
    9363,   9366,   9368,   9371,   9374,   9377,   9380,   9383,
    9385,   9388,   9391,   9394,   9396,   9399,   9402,   9404,
    9407,   9410,   9412,   9415,   9418,   9420,   9423,   9425,
    9428,   9430,   9433,   9435,   9438,   9440,   9443,   9445,
    9448,   9450,   9453,   9455,   9457,   9460,   9462,   9464,
    9467,   9469,   9471,   9474,   9476,   9478,   9480,   9483,
    9485,   9487,   9489,   9492,   9494,   9496,   9498,   9500,
    9502,   9504,   9507,   9509,   9511,   9513,   9515,   9517,
    9519,   9521,   9523,   9525,   9527,   9529,   9531,   9533,
    9535,   9537,   9539,   9541,   9543,   9545,   9547,   9548,
    9550,   9552,   9554,   9556,   9558,   9559,   9561,   9563,
    9565,   9567,   9568,   9570,   9572,   9574,   9575,   9577,
    9579,   9581,   9582,   9584,   9586,   9587,   9589,   9591,
    9592,   9594,   9595,   9597,   9599,   9600,   9602,   9603,
    9605,   9607,   9608,   9610,   9611,   9613,   9614,   9616,
    9617,   9619,   9620,   9622,   9623,   9625,   9626,   9628,
    9629,   9630,   9632,   9633,   9635,   9636,   9637,   9639,
    9640,   9642,   9643,   9644,   9646,   9647,   9648,   9650,
    9651,   9652,   9653,   9655,   9656,   9657,   9659,   9660,
    9661,   9662,   9664,   9665,   9666,   9667,   9668,   9670,
    9671,   9672,   9673,   9674,   9676,   9677,   9678,   9679,
    9680,   9681,   9683,   9684,   9685,   9686,   9687,   9688,
    9689,   9690,   9691,   9692,   9694,   9695,   9696,   9697,
    9698,   9699,   9700,   9701,   9702,   9703,   9704,   9705,
    9706,   9707,   9708,   9709,   9710,   9711,   9712,   9713,
    9714,   9715,   9716,   9717,   9718,   9718,   9719,   9720,
    9721,   9722,   9723,   9724,   9725,   9726,   9727,   9728,
    9728,   9729,   9730,   9731,   9732,   9733,   9734,   9734,
    9735,   9736,   9737,   9738,   9739,   9739,   9740,   9741,
    9742,   9743,   9743,   9744,   9745,   9746,   9747,   9747,
    9748,   9749,   9750,   9750,   9751,   9752,   9753,   9753,
    9754,   9755,   9755,   9756,   9757,   9758,   9758,   9759,
    9760,   9760,   9761,   9762,   9762,   9763,   9764,   9765,
    9765,   9766,   9767,   9767,   9768,   9768,   9769,   9770,
    9770,   9771,   9772,   9772,   9773,   9774,   9774,   9775,
    9775,   9776,   9777,   9777,   9778,   9778,   9779,   9780,
    9780,   9781,   9781,   9782,   9782,   9783,   9784,   9784,
    9785,   9785,   9786,   9786,   9787,   9787,   9788,   9789,
    9789,   9790,   9790,   9791,   9791,   9792,   9792,   9793,
    9793,   9794,   9794,   9795,   9795,   9796,   9796,   9797,
    9797,   9798,   9798,   9799,   9799,   9800,   9800,   9801,
    9801,   9801,   9802,   9802,   9803,   9803,   9804,   9804,
    9805,   9805,   9806,   9806,   9806,   9807,   9807,   9808,
    9808,   9809,   9809,   9809,   9810,   9810,   9811,   9811,
    9811,   9812,   9812,   9813,   9813,   9813,   9814,   9814,
    9815,   9815,   9815,   9816,   9816,   9816,   9817,   9817,
    9818,   9818,   9818,   9819,   9819,   9819,   9820,   9820,
    9821,   9821,   9821,   9822,   9822,   9822,   9823,   9823,
    9823,   9824,   9824,   9824,   9825,   9825,   9825,   9826
};

endmodule
