--
--Written by GowinSynthesis
--Tool Version "V1.9.9.02"
--Wed May  1 23:05:07 2024

--Source file index table:
--file0 "\C:/Users/stefa/Documents/tang_nano_20k_c64_dev/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/Users/stefa/Documents/tang_nano_20k_c64_dev/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.9.02_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
PQ3giQmdEdHWU1PZx7Vc3NrbTnuufNtoiB1jJOWXM8eFeGbFHgCi5lddFIkGocNZxelVsAdLZGSF
5oz63FzkrUCKlPc4zHpZ7P1HABEAsE8hMRBMJHEnvScNLHqDj1dUeANIliYNMK/s/YNy+VLgC40A
EI5tSYcgkCP7EWy1FCrEfl9J7I+hyYIsOKpE2qLZ+wwYGSYw/yqWL23V9rHNXsTF+GNy8WT4cYXy
7aiN3fIelQlE4a3E4FOZYX0o3GF7B/7d85J+zZ5md2T78l8phzGwseKRDDsAOoMYzQhOsQj/OBlK
I5gO2mS0b4hDOp6GXGokenjHGBLD6L9YYuGbww==

`protect encoding=(enctype="base64", line_length=76, bytes=11296)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
bdEevXnuRgmLERFLG6LW0SlYpyJgwfV1sUVlayc7NMy45xZGs+TJADmo+FuzehX9PMIpeVZTnF8v
t8X6EVpaJx62mOE2gCHIlR/L12d7Tt+4B8ohYTAeBNMUZpI98sdMaWIk6qEa5z9/xR3WecNbsVez
nm0umJANILznO4urTClObcVVgZAaimEKHaTGe4NtitysP7brTkAHwKDL1z7zQg1DfjWaoW6tH8fr
XpejXjsEEGM0+X/dSC9aQo0BLtGFosPwKZUO09xKDWE/o6eNoGlIbcJWm6pNxtopOurvg6KoVPEH
i7AK6IhUM4rYYT+H+a3Wz/mhIfPqI7HBnRP0uVN2PRwLetGEUbR1y4Y0/PAqgwgCWULlIcW+LaKy
X6PPBFMA6U6MoFxcujFROLIjAaLO2qpN4n2j+Md/1QPJbUDv1ld/UKrHeoqAwboaWf5ttzKOLfeX
i1xQE2wAKyg4NwKqFJRtC2dUBcS+IeNU4KJ3oAc+HjooBOG90EYNdRxkLwEoU1ek7GrR/i+RgEWN
SyfYakuWVtdq+6PEEJLzbgysM2vlGTF6p3Whmt61LnCmDUYmDabhKTRROg4qyAnr7xXBCxNDazjK
9m1NI9YhSL6QHFl5OIfjVVwqP9tX00so7dZKjGvJaVjnmdfus+gpQPsltBpkTti9/ZEICIoTwz07
ahmq9bV0W/1fmqCw9P0L+s9ZUVCjhXvAJnuF1Tj9ClMMvBgi841A6mOVcKc88IVu1p2e1lZts9d7
nt9srJCw9MCENUSr9fp7y8IJb9i/IAQK3zA32rU3m9ZkuR/uEut3WnbRKTLC2gRGjGNsk2FE7JP+
+8h4GREK0SYfZ9qzG9H0X+I0iSOnDjavQZJSTJjLoimqmWXEqmJofhStzb4MEOsa0PnwOZ3PCL1K
LBqg/BevySS5CZ5RhEnOfXfhXjIDA0faBIMmwaUrYdlx3y/jvRLtN+3cRGgcIiobroQunayYBHIY
IAAZWggM++AUYshvpjAB54/iopoS9eWty77ectyF3XY4yy539u5nBbwJAOu+MxVrzntu+IW7lWub
KKRvhKvK3yzACWF/W29Xc594xlMk4q41GyBPRU0YPZxRcS0O1arHgLlGE0Afj8Zvhwxfymq/bB1Q
dbZlVlFIAMNJCA/CTZlYfXwaUEMZcJruaUJJ+3Muh0njHgvvcvhkB2TyPIDkv9WhHkREfmcmbVJl
CgiG+AwfZ2rUwpIFgpXjLD33XB1rL9T6eEvqNbnwZhPZZ40wzRD43bIf9Sb1gFo9B1Tq5faWvdTa
Wsg0vfm+Vxa2pcg4S3o0tAEn0Mrk6GcVazWSdRZxJhizBuL86Ia600bLEhhqZMLEu2lgmzhhXGIe
L+iLIxE5HJ8nmjMbtiUGH76NAgfpGxEoLx08JJcpaRS+cON79HueON8KnuLReKvNERbeKrss0e5g
z6pUyu+GT2iSgWpoPzJKlQVTrYk/qZ+rX5VDMFrFAGvRGU1KeHSjbSqGYtg9KuJkvvPFpa2S0ubc
UyOLdrC4I5zBtWiKW7sed3JOh0oZvSiPLzt1PNh0QDTeM5a/RbdsWuH55WfsZXWn8Ttj6Q8TB+yX
9w291jNtLXO2YDqTslJ/uRXAOeArBrvzU0pEhOLVaoMefbdE0lQCgrkmhPw6KYl1G8R5HdCt4VYv
AziaFGSJX1+yUETMwOXVC0xxHZzb5R0XZj/LOrTL6X5iEqrGK+/yxtnZo+aJz6sY6qUKRovuOb0n
FkmL0aiRjB7FJ1WAhiBftMHExTBkDjcQdBb5qqRGpTmodigVt3NFVCHw5B7PzyxiHw//nm38O9OY
iL7RydzpPRbLyIcOOn16riSH/kf6rocuqF5HJJwAF92eXQmRpQu1oTTJZ6G2jkvG3+MOblGkUgzN
qoqKn1a6w6byJe6Z7zmciBFvpgea3IchMVfMStCF1HKqTiFCBCCgxSm5WfVOmBKuGRFkk6ontwUu
lNidKcFs9HNEZBBvZgNxJtHJoo+ujinfcYQ6zGR05GQHgJfyNAwpsb6V9F83hRoDBHAuBuCW35vy
0mW9CsQy+DcCQuA5QExQPmD/8EzYWnHDU6TwQWSLdXAiiNSsZaQrNuZf0xbQOoRlgWZdiOtIHnh9
+NSoGOW6LaVmefP83q+rgypF1/kQyRSpfr30ijIgw1h5kFapJepTt5erCAGWYpIccY/6PBQKoCMm
zBfh7kndUbvdtvb3HcKGd4ufBT7dfyAA2EI5buCzTPM68HFtbmc6pzpL18LNRzhnnni7B8QaCMiv
tky/611N8wno6xMsT0ckFCqDk1q4s8NFdPe6J+sF4wjjpTP+RLgGJjrU7yrv4DhpEr4sMUnsLtyt
m+6kMwsLvAPA6+YHfQLU7FpP2t0mBzsQ/WYP+7ZR9VpxgTLT21Zj3uPlwuJIXwc49hxI5v4cDnyy
yfMv+1T5OV5RBn4VE14lvFYB68+hRQL8gg5W9wLfad6UfZjkNz3nru3r6E50Bm/W0HlsrzMJQrCu
A69H7MiLrfsVmXkNNjVFQeXWmiJKzGXo6/ijFYCqSu8ZC6VK67XO8n81unO/XKRVYIF5ubo1zyQ5
d0cE4ai0OBwMDMCSjrPAuIoUhJqCmrv25MrEVyS2Cr4KInsFyIAHgdtBIRaTL4d2oevvXpZ40nm8
fPfmgqHZ6byqihWHTWaAvDZzQ6mJ8/WFTspDB1ucQjgqdQEyoU2vGvJVP/EjGN1UWn4R1DQXHHrv
0xKJmk2h+HU5XCu+HyI1EiSAn5a8p8XZ+DV6NNdsUPZ8bR2rNQ1hZve5xEedM61vytxK0QNOt8zk
0SO0DRW7+lahZEDhoHJ+ILHOUne23inGpFY9w7dnjbL8Dat7yN5UK6wN5Ka4GEmfYM8jhjwHkczz
3yTqzXzN7tUj+g2hIr+Hrt20aKkIq4XekEa/ELcP5RfJzMaWW6cajsl3bB+rEdHzZPP+be3gRhwJ
XHxiQt2hFN9kG2TUEzoUeozl3GOD8ItVOqMR0Df22870Pg5YCv+5s7D7Vda5wAjmo5c95Pdmn2a8
oelX7w6JJfEhvSsjxoed+XO9NdKc5l6P0r/pk8FekgjUTUUGm4+TkYVA8neiF4YBk0Y+aK3NNYYD
eWDUdp36bpaoLoncwdPXbi9dhrgtB96oJU7UkTDGo3Uj1zSahw023SP+VaVLTb1+r8CEhaiovtPA
bRQE2zjQaBV8S7U8WQaYky9Fhyk96z9Tt4JReHuJQDLqwFRsJEMOqt1ohOyM+a9kKLn8UEqqm4hy
H5NxSp8Fa8jQ8yatt39axvMt0lF4qdRkuhjB61NUqLShA9zT33eESEoCnx8ERn/onUAuDgd0BrI8
o7PBfE1EPd3fXAryEaqleHrkXjutnkuyLpnvYERsdHkXKxc0ZhC4X6hXyZjTJJgM9zLCoGWP6U3s
9PJPsjXd1r4phNvDYune1Z+kDDxLf2I8ep+mBOKKBIFaPxMynFbzmlfl23R753RcVblsjvqeZwZO
jnhedsEpKKrixpJiBn7uJhBOcrh8gjgckZAEbt3oxvn99BAeGU9l++LbZXai6edE/bhOq/j1X5Lx
BYVia3sHNUGrDDi4k8YbKgJa5RJTM0tcmp1ZqMhZEohKKBy2qa7lLNrvljtQN9vNkYEJq7Y0thkS
/4Z1ooijfZPj1kIrhwj/LCR9ZGx44JiBd3V8QxU3oUpBFoNrdvZMJIoQsC4WA8iRRu0Td2p6WCpF
2iLk0B8F+F+KiY4XuVccj8t4OLy8q1CC/1CpWoCFAF0g2hPpdpRlBx4RDVycwoUVuwmlHiaBFD6/
Smw6ybETOTHAtXUcXICMmh5k6wunRhJFPw92GIAZnk52ye7GxbC6MjyCEZaMPoIZAI6OtI6dvr90
33CBFoAI4kUnk5IR5XGX84FikhGzwimm0PfojM12Q+dxWAxEDHN0dbh89mkHZ333PQwO9PYTBZLv
bO8Jtsukejy8JsU//5Cu+ADUTu7sh2hYUWzI9gcUbpQIgtEAwYL9plTYFxeN65QMlm2LLx6eza+P
R9xschYkfDJFbSWmeLA/6PWUfoJWwiUtCjddm05+bdcKdfbKb2AmUOoZlhT6PR1bUlwxUYIhIgPO
qLLLfmzjqvO4qmZO3lKSho2SYnprfw4GWSpQazxZtvFD84MJ7rhd5zlzKLteWesdiPO1TmDVLEuG
2P0fdq9g8YT+4pf9uKD+z7v6EL3vGsC91WZIYY0+7IKjp/Vh/g1umrefyivRumO6zkFhYsa3iN4L
EaUztub3OgiDcL3dvPnWUxwvUjgJHEsO+PCT5bxnsv+wEJTS4h/ZDjBmp3eysbFnjUpBoMPzJOHp
GJAkZLTVJs0JMhoq1MVKip2ZnQaATcA+3h3SH9GdEjGOW6G21iX+PjKFSFwLSPj9V6crdDrP00Ll
wzr9+XPRoFpuh7g1gzXtHkLJ/tRrW7YubOd3cGh9tUU48CriYLM5xw8Y2f/Klgz5nX0kNY89CdtI
iQjv9JBHJYjbhBXVByCUmUUCogjXXZk2cU4bMtJlIeBgqJGGiDla8mIzHwE6aYTmdilj9dlgxtDG
XX+4rtFFAh5capynfGJsgqOwgVPTWWWZJldliUPrpRCeY4jHeLACmLFP/IggqcVv2qcKjrzL3Xdm
LaFpjxWQY/+PHLZPeTGyXlf4qAP+pnpaumUM/mitmxmVK+VE5L134+I4rI7Pqalb4yADlhcru8HR
kkivjnHbmOj4CM80F+LUEb/goE+I2u9iKyNrZr9gmtX2ulj9Ua5v06j9YclUOimJKCy5s8EmZkyM
wZxgDexhxnRwUURPfkWQ7fQ0nZdcNt2Czi8NeCrqkgTrJ6eiD+uVWF0XHR+AFLXIA/cOqKXXYiMa
+pB78iLukLka7DmmyeV9ZwC4H8d4DdJKokGfU2mgZBXUMjNgoxPWlOOpyOMU/ELNgz8mICfpFwnK
u0btS1Ij2xAdBy0844Y+m8W41qwExdXoJT+41d6AFWyiFAFSPyF4OGhvfhzfwPuUWImx6ZWk6dFC
bOstNmh69dwwz3GkuphwJOKPzJTWlGBjfq2abLbbQN99fC4hk+vj6OeDmdAUrVnof/ctR8ZOdUFH
MyH1Lufrgcfy2/N7NU4KxY8nweG01weJUoi1cyt5OhkWvNMM1NkxlH4n0DpHqlBJIMhxSqg+1VZC
AGtNOpIDIaaLx4HhXTHjCgYfd5/hMVLWf4GHJBQwgRgzwhhaBaViDG5SNczoz2uI+j2ACp/1s++V
+qNqYFDH0AYDmC0GKyaYq26kIvdQehjnf9Shkoa0RxGdqiqzGS3SCS5vtHjyTGS6DWO/PPfbLkDL
xXHGCV/9DA5iY2hWjpqno4oVEt4E8L3cUJjaVtVFbD26GZlbr4nk6JdDTfk6ktZNbxFVccaJrLcE
x/uF2QYwoYmHiN+tLkcJC5f4919rcPLavfSDpKDzHTPU7k4VVOMx1YFPqgmOqk1EataguM6r4kP9
sQqvcMW0sOPjh8+92w0Kt0BHVkttSIvu5Sr5qAwbLtmBxIYzxtBu/83avW0MtIsm5AL+j3zSkBMa
b1olbBKWvk4SPAIL2b892ycbKn94RAvTNtCZ0DnWhTrQwvBcwtTxKKVNhNRPrr+/Nqi0yU/6GJkd
7M5ybz1H1VZqCbPigKCJ3q011h2BIkNqGt99111XY9UpKxNTXw/4NbxSM5DgMslhgq9wi9aNMfmA
aIHwslDoULU3hhroCW9OL0vlN/k4WGMI/mQPT2Hy2FtSY4HbebvCLxPTp9UQl+9KEGXyzrjaE5qV
ILj+HGYSWfNzSTzZalzzql1zYc6uR3RyK1MngmEP2tzeKQpuuEjqDp1YLnGyDJS9lSaKTN+4L5QZ
N+S8vfarFmBdia7zeB24XImjYSGDzUpLDFpcYmgIPBC2C3E6RI+hy/z9dOrbLgiZdOUtKt3UirI+
FHPH1kROG9WBa7Jm2nHYM+3ZvCMhg/sp7uvo6CPyn3vwc92jmwbN/I4asLdKBt5YAl4JAz1J0cEM
St9tUzAqNv9UkoH6/5h97F5pQEoO8xoIgduYm1f9VNUKZnnvNrxawWMPbJKbhN3Hm8LwYizDW+Ak
rFg1vPxcUcMQKIFF1+UyGxhxKDEBiO17HTtNqTzl5szunVSKHT9rfudamuOxrEyjdtB15TXS8RRA
rtelWnmYTSv1ofy6kUypr/xR7EWD+8S9EJ2sSFksfh4vM4y3lAvTX7PD8jKHSac8Mri1ThDKCjb5
vmIAMOn+CMFBWqLBLvY8LFpcJLYLP/fgKzDGTLoHBaNTixNx8ccFc/BDFRsVkGetkrRyvZFu7wHV
yodOTLG4JUChFkmZWRwgWz1aXiJ5vmceNW17aYr8Fo4TKPH59nLEn01Ij4UVxw/y7+TsArwNxRtS
Dmnwnd45siJ6wBhTw/LR5DL4k12cQKG1NiuKYAKfqp2aC1cXuIOQQdlB9mbv5wSNV/+UNHWiH7HU
eIuCkm/mnaKLIQKY/MsCTM8xIxIm27yk+hlDmy85vaL3pz+LjP5RNdCBnjyDFcoHDcoCoDBU/207
6CZNWLV+ABgQEfvvo5wenClE99SzgRBo93zi8tNxQ6CK1JWE27N7O+U4c4lSuvdMyQ0ie7MXkbEy
NKBuMgMPUZCUXBiMqQy9hTRSM/ZZnY81Lwunj3xJGFSsNfxF6O3HOButzuZNIK9Pr9YzADYEHKiu
/aiWzk5MqN97xKT20pIuVcKvWFcf417+H31JpZUo7e0JN3Pryq2jOqODf8bQvIFHDbpWwyWPwrnI
kkbR0co8vMu1SwPDgAvuVe+U/yIlhnnUIOoy9rrwle+gbw4IQ0UXqXqMaVbWqfAxGpngVaPDHqrK
AKKBGdR+3fZTbb9zLmRBqHN0qhEmFBGx1EZYJha/yO4ZFU3u2rvl4zRDm1yUA1+kkR7dsJTOmgP5
MUaLUvmGqHePCcjhiX+WZKXrs/5eFJ0BeJhaGw1dqe1ILLdSo5kHgu1JTuO4BGipCfUzff6K8ovv
3y/J0dWLU/6KEldBhZXYiRMkhzNYZ9rsfFVRIFzdbzbhOwjc2S/Xn84ABXTStlkeZfH0GT7Lwqqg
dIade1DC2g42pdUiw7otX2vmBZANyEkMtjbXpOan+UYpw3bMf3NNfYgBt6edadwqhe4dOUhlpeCB
bD0MinEYUaR6MsKBry0lEXRij0cy6zETv3509LC3q3P4nBoDC5Uwi4cC9zQaRB8Dk/1JQvkGmkFU
suOaMp8h7ggf28RBAtjVu8sSBTFEFaCc5DPeqjbVhEiqFVMKtsDsylPP0M7wr+Dm0bRsg+AxNraL
l7CQj8nZrKYXDFo93mOvR8twfUjAtjBy3QSrVb+Ha6Ej5CBTs2vqbDBIJDZKOUWl9Ig8bBG7+xOV
NHuoxlbE0W1DJYd6ba1HufDex/avU1n7hs2wlDdAgRYUVOsCO4T0mW1oaZ6T5Hkxs7HUMQIZTamI
iZ9KgRnPhhRgfQ7B0bf1Bw9UaXRlPDxDfb6QX25L2MZbRsjBD4YoU7riAnLX4IkBSy6vTfNj3+86
C4lx5NSKLWEtTUj6l5nC0Pj/2bhEbhWh63rxkb1mgSfB4CPUBrnHiHicUaTtobOzSxb3VXvZ+6/b
IrYKCDMBBiVvm0hbRJ2T0KTGdnAJEPBw58gw/K2Jwx6VCiM4zGESTBW/zSD7CMq0a7Vt6V6CpsEd
mn04kyD3CcxXIvNnG1NRfBwi30b7PsBcEWMcnIlMwTJflsofe61Zqnddp7nnPmJIBmNr0Er/MhNo
RrptxYPWqjNFz6cuxdbP7UC6mpB9NlLWidPFvLd2zA3eQAnxXxEJ1wQ/RmHYdznnHoHDnS1tyUyP
/uiPHvAKoxQp6244A70moLcAbmvemokFY7lyhK52/4yQ2+898f5UPF0iutVlhdOhd0ZzYn4mAXB9
VDQe2nk1+igkV8fu3EeLCxa2aMi+jVvu/BUyaZWtwnj/2TViVnxo5ptW1al4G8d2VRG2os4nq/wV
fIDoJmoIWf4WxcFjhffgIyhfrlgA7YIh3bn2+ezvbq1y4CpuZIHoqGguLLPL0sAngBEIkZsF8hsp
f9jNhaqqfZaYRqLD0V01VPIA/a07sSEHppUk4L7IRSFEHf10yX7Rufav/guw1emqWZgPVTr7v/qA
nndKZl+QPl2Rf+/TaOcawgid6Yvt6yZIjVfc0gVWNkQfhbe9XI/yMBTZA1iZlBsFICi6ROgx0kSv
VA+waAEEpG6NZHp3b24gNQs5L6asH9cbDWncBd6IMIo2P3riOTTtbKD9v2cUMztY77izdE5DA1DH
8rQuI/9J5aHfa0jdXw96E0oELUHo/Y2CmB7OZGcSaE3UJNW5nQx09IKOqx8RShP2rTs8OYKw0hNo
njALAeJHkNoIpzzS/sCF+H7OJUHfIXxYXqbTAxPOxN3eyPbph4hgtJzs7lGInZTBY53/9McoLn86
x84uzyhmk8yQ9t3E3hk64sQWfICiqHaQ0/+XaACZ4jp+fzZZWe9noTKhUIu4VHnCN3ZvCKQ2CnP7
Ieu1AGr818yr4uOZ7A6HO67U19sNMXInPwbudrqyrvAR3jVH8a8Qfgnv2ctH9vDeaxXcxROT3X8e
z1C8WqOS1c4Z8JpROeDS9EAkGYiuOa/C+uVc4ajLllo5HPTXJWldVWNJ110MuVAagUX27O1adYgm
DggGMyPaGsC9P991FPamAGSFVLBMgBiv0ohYgaSVQM61mkEMro2sqaAdDJebnWgy7NWgvg0fTuWZ
+boxV89NqDB9A5PEFIqM/2uxLbcplsc+RlUu3dNL5as9OWf2Bjqar+Kr7chsmxjRTFWIxMuXEngg
4hsXAinIqoE9hDBpTBkU1G+IOkGzMZ0D/uISRwWWCGdYA74WTU/LJmyQ6unQyIfoyK0gUwT1kVA7
v7el+K7hrHpDtJljx25EYFaAGQ5HVBAYp6GrT/zcV+d30dv8H8DaNDbJFESskfubaOZaFxTMuqmk
U2aPyCY3RUFQoEvFlGcv39pDJzcB/UU0Wr8yxEJYyNKcpv12ihBWzf5J8uAPDv8GopYy008uy+6n
dL8yFRqo7IL31nETihqjmR/+zzQ33MJZiV6ntwhaWm/rxjoQ5mlYMD1L7UUl+agBx3GQ3897UeuY
16uSRRaZH1skr44WIPm6byEM3mbndz/jNeHhhvwVDlglwgw+ZyqnKkJniCU0I3PhYVuiGuvFnA6h
pe0GXiMXphrWXokLxqiWY+7elSWyrGTMCmHVfsj8qsYXrmm1eZnZVLCzgB//VN/ws/cXJv43Qt7H
UwrWbv+RQVGw9dv9vclMR6zNk9uvGLFiOa8oRh577hcCAjG7he+XGr5kKq7J8O/bLi/pzBjGA7uu
Z/bds09DrPGNF/P8cZAWCZrFUIn5KURfOsEpxjYwDaMTsLrqHasofJbixc5T2mCfaGTwPZiz2FTF
1CSdS860GJQn4Fs8bfi4WC7n7tTRRsUwQwDiatMu5U6Uen19RsWda9pW41n6XPKRkeGzUfBOtbXn
i4vSn3HQHHsgf7wT9Ml94faztONdloajyyjSA/mQhEiHx93py9JlUSGU8HuPWIAc8b5PnmbmR+QS
n/RuP5GOHGwyGKcTsLxSPCM0uqB2hIvoBNYBwEA0DxEDNMdLcC/Ajs4z3AI5oBCklrASZ+fGmPYU
BC0aMrmtgypH6xuqrRoVXquM/82Ai58pHoaIXqDntjyJyeiMOCC3dQGM4YCw6ZpQwMsDOM3WusO8
A7autenA1b1kDjuW3FYKZluarNTQ7lHEcFm+4TpIWGSXo6xQ9ZM77MnX+FEgVaTUyiFTMydlIWKx
2zFaK0vaNhN0/Sfio7jyGhUuPCHFon+LLTxLtf6EeARb2e186gEQ0KSV0UxFSZvZoPO2q997RK//
pkxbmE3yVCRiEhXIraI/kQPxtbPWKFx+qENRQY342qSV758qYh09bLLlwf08HdtgFhiLv0vzjSRD
pHQRfFIIu9VyyBfYID5eZ1ix3tUt/o/SPA6UC4bwU8eI24SVvxay7HKr+QAVg5nEUqsPGKRbvS0X
33d7NCEf4McD2Ah64PLeWO5+PJzAEXhAvoKALteygpDNrGZV80KaHAqEOsz2ZGPr9MtIyvyiFN07
XTG/bIFsUPDTKKzN4/em4m32bM9Ea9Cl1J0DDecibB8zyAtmO7tlecXux6SOtCA9jNObpqo9KnsX
W45t7JKnfdZlPnW/Uy1T4HcpVv0rIy1rk8eDdq0/j2hzhdfa0NfHpF4Yvg7J6ukNR+DuM1gRBkFG
uBaYcOF+KJXs21g0FKw8oZndBreLmcUEldVZuH1ixUlzoVPbK1DUnc2Fcivx6i0/OCMON4SfSFBk
F7FkWYNM9PRAyGaJUlqJuwgG1V2Qyk6SVOajPOS5Tg9dV2XpIiG5payqI3/Bq4/oIHV9bazPDZKS
/GbAKrnkJMoSD9/wJSkumeWs8sVtudAbgz4U/nHQPwzkTMOpkprs3xV2/p1FFLjkjWhNilwetavs
HplUs4rhP/NnrmwuC+DF7kKRUoRppiF5n9fiNMV/7O+o+fHASoxZ9PMCQGvSMsfXT1CgsCF8hH5g
KkPVXzMVTvK8GvBPrbH9tKwcuBu89fXU7IoJ4EfmXL5h0ls3U1GZHLtECPxwquKbT5iXve+rTHMs
TUmy3cwTeGvBhT2VRB2RfYRNy5ZtKRbLqBAEbaZcB+6w5H3KJM6fEO6o3GTgHDZnQRRdQiWP6XBx
pJFcT9KDMDptPKlqL9lfSXUVWyfKJth+RTph3q9YWtXQWasgo2Nycn033kR9bnwJQAm6q5NNAAyv
U270RUE/OchcxdAfOSmsxXTDsrbXA4s0kbg2ObFJnm2RqLo/0TxdiqlvRkcKwtvTj3Tm9wAPWOr0
fZs0RCRBdlZPhnExaphvAmVTJ+8PjdmcxlvHtqZRmQtd7cYBRmNWJJUuKbS453tn+gaYr3z23VV6
SdD2A2F7+Q9FEGRoRSap121q3Q0XpmnjSNoFfVZpDA7lvxWMfSBlrZcK0hO8oDiR5VS0zG1YbWBZ
uehm1t0/BAYymKsJRhGgslIy0AmgftqUrhSMfOtnHQpUEM3yJD44JxmfFkD1JCr6RRgI5abEfk7k
jWo1akZoMlw/aQwzm9S4S5bQNsirzEFtvYkCvEsyx4uRJCVJ8agd+abKYZ1HCgXlDBd0n/PoJn5l
qxSoo21xRzPNi7Yk09r7GsKG5Qe4aHtFMeJIpd5fDi5RQT2PN4RQQt4d7Z2+lYkamEjxnVhRd88Y
d1gtByvlcKNOSd/0/FDQgPdh7aFZRPlDZElIO41oGu11+br7T0BnlpIEth38SWU6c/esoveNnNkM
gD1ned45zu44pCCxTyBQG0WZf9cXiXUlD21Nd0tBfdRTStSDh4e5vasOtNRftBoTK6YkmlI35eRC
ujVTugOwDR3k46AGMoxIG6LVKfxhiIdKYf6cIw9nbmPXbigJv6RASIxz3Ru8teSgZ6rCn6WwGxM9
95p0n/wkRo343cOrIfoWXC76lHuzUWQ9IXTSIqSvqQR5E7m+KIurimmbJHN2IUVGR7smhf5s/ntD
h9fOFTRVXNCqO//LACjlNoUuYNWQBFz9eenpPqq8RDZQx3cSVEu7Ry9IQ1Rnjpb5eH7hG1ENDp36
U9xBQ6qvZ9mSmlRQuzWHyyn+Fi5m2neoUYnlx4uQiyNwOWPZXse9TqqzEQW7onUoJ9lizNjk2X7T
dNVHq6/qd+tkTfgEdIradv+90GkSxCrBUeVQxO2NKFUIL5lFqWYrQkgA2v+PVr017AmM58JDan64
Es23f/G0S+XFPnO0wYGYtpTE7vxmaI/c4NQ2Xpqa7DZ7TdQRZdxHxGd5WzO8b/6yYuADzDuhlPLP
z8QQ8eKnAQD/dmsNCX7jITPu2F9T8VBkhG7F4ZzYq6Qpe8+L/xgoMmEq0v+CZCQIytfa8A7sr/Io
2K0o4psLk9fB7h5wH953Nh6dRJZjYtn8GAXEepexHczAneo8a60OjmkOUsBZqUhjo+fuMrBjH5/Y
QwsyAe171PM64krJ+71vu/8PrQLAkVdwVFJ2dEx1yL6wC9P4hZEK5X1gONjaWGqcNmdsKBKbHIEf
EgJH1xT1gy6u3L2TRBONiaAomzQKOWhnXyTvEU+EC+nA5yTbplzGAol3I3q7C+CEt+gOhKIueLP1
qJq5ZUgTMXW36V3kTPE6zJzYxE7E/ePMEiFzqQ5w6Z9NW6ZU5lFDz5zwYmcGcVIBUj8cDCDXi/bN
uQR/o28GIcJ4TJpx85RvTnMRxxSLOgTAkXFEV8TWhSQm+TYobDO9gLxpuWROKWnuGoFqdCnr62BQ
1KKqbh0O9bvd7l9TLXn+1eEktGSzzmx6uIvsMtrUpA/SR5TB+C7pqFgy9K2D/21e/8o8cMI+pWA3
YpEJHdN7IoBY0wpXsYx2njyUkVbHe/SlAiQcrmcE6xfBG7nl0w/WfRquqBEREGJ1jTMnMnwxV8Ix
UC/XvSJwZ5ieqoR1lRlDTBmZ/YVeRmyo7bVAiejSJ75eZh9s6oFRCtSW0cdn8NKhGcqOGGIfbETQ
BJ4XZ2Z8hb/QaJIrK43g8bMeFlsaVGTZpUC8vvZkaSR60GZDYI97q2JybKY7pFzu0aP6US/53ngE
svLNO+5+ohrLG5EfK4ZQ1yb48nQ/AAKZ+hVaa+bj9+nGeSA6tHa9qFIvBz3xNnKcgVFj5Cc5CYPd
5u6P0jTM678I48qeypFtxJlgdJpCNZx8MF6bG+Q2chsplQJWmLpWvaxDjWB8IGLED1orr4AMjNR3
EnqW4ZubZvyLAyADDhBR2dH9yMtfxJCewGX5PfvGzB/Pf6moIRTqra/0tKnF1QHbQUaTqQ+bhWis
Y3GNDNUO3Bl843E2qSrtNUCtcpuTQvFlGovPykzSu9tBdhp8e43ikp3sqdRLcQgdbrS5it6xKKir
S5WS1nmNkslnE2jUOmwLe77pfOCoNJtGGWa+EYz+ekBY1vAmnwiKAk9gm32bIDE34wEZT+QcfxYb
5codhSmO0m7id86kGxltY16UNCc1OTeWCluBiR0jY+XP99VF/hl/i960EN/zuOlyLZ7jw/p5FAlq
jQu/b2eaWsFG8rRbJsg/1MDsGEoMCgL4EBRALIwfibBFEMppRtbD4GLxybb8bmu7J5NU+Da+Jl8U
hWJ4j79izaPg0i5En2/XPliPbu5X6RQwMfEMtyyHpcIOH8vjTZbbN79QtEOoSeUDVVOOR2lPay7A
kLy6stx9lOHi/Ow4qCav1HuUr+yLL756TNVyHuBvPPAJ3Wgag1R1u0UhU7DbQMMKKZRBXcQmEnMw
41WZpFjKgsJ/WkXkzZWgvUdNJBAssoAzH8AiK93ouP1J1+dM8v6vQGxQWdKoPWNekgfqym3uuL/Q
f5FJjqc2JGTlB4Nd0YDOn+JgrjwN4GZcMPvKb027sgU6nFos575Sv4lL4cBQTAStg0YB8DUPKNtC
cNR9wJNOYl8J4ak+O7hx7myMMz1RfiFyiXbT+3qTvDRvIVyGuHrWi5uXC/PQLMox1xs68jIwlxdl
d3Q+RBROyryjO+A+APuqFyzgBgx+MR12OJ74x1Iq4GVs5PIbXk6/IWKLP8nCVescpG90JI/H6MvW
v6E1s5XygwbAHMsCl4fok2X08PFs+tLVYQnsRTDi0ttN6AH16/QJQ6BJPCnuQ6eBbfUVe2Yxhbvv
YnY/ZJbI+/t3NLa0tQwmN6GgZg84IZvCL4YrObFyClTIn+14k+IqN/gRT0mQI9PmP0K5IqKcT6Mb
YOz3vSn4GPzpr/MYt6arx68xD2mgrMlBKQKQfpSXNlV/uU+6lMmFnLbP5eww59pqUnXMx9fXjdvW
Id9WKffIQLB7UWsaF0qkYzOGuGtUOjGdDv8zktG60Cf+ErAByKvlBh5CXJw+/n6QaBpnPs0xeU7P
zAWcglHi35XCuvhm8AQrc/tSgbNKccGJck2Q7aWvUeZ9Sm/qOyQynuoGcO6/LPaxkvn5jppEvVUU
9aTf/SDDNBvnCS2cHuxvW7M0R6Kn8vNmDF7sNPp9G5Tq746TGD8v6VyfT0jRKtxlqjrQz0l+8B8g
8HZ/kZWNfn7vcbQ/AGXFKBaS2dr9tcquj/RTcFjgrU6ZiQKjDDfaYooi6hkLY2P9RoOna/INtaCK
SVNIBzzb/dHl4YEGy/xEOq3o6Px3b/sJYThohEcGqiDPJTa74iXB1moXfabqaihwDXqJ4xBpKWOQ
qkjxww/c8dJLFjuFPNrAKCKJk+EinVqDY030SMworWdy7VDqlv2jzBZpwZhQNrcanaIIcxB+j8d5
/1EYE3+LB+F+0xH8pvQq068984Ipfm4oIthiFzYy49XBo2jm/5Lh6dwhtJ0VEZr62t9ayCdPxYwA
KW1IpSpRa1iMGJk+8ZUeBTtxuFMAcDtEQTTvP0LyFU6AtI5XoKDDh4BrrPjusrPxrlEZrX68EwKL
EuRd+HNI125jPLdk7Oz4cDG6MTO41O5hNW/rRvM7tvMSJhmDb71RLepYuYfF0DmSfSHYAUz6gjeC
4+3M6Zuivv+2cKG5NnW8QRDBvfM5aejXGvCrkoE7NPs8wqDpDMaHUmtL7r6TODTM8Zm+FTYvVrDJ
xg5JJxsveqOrMB18qVLcE2IuJh1dKfo7sJFPQ1JmwSK3Q/+f+AfsIXkqI2MBf+xqGyg6DHcAdWYp
maTaUVL+7eKJ43qasA4AKKRe7vGQ8k4ByYUy0RePuaKXxaZECRdy80xVwCYd5MoHGTBeWQxiVep9
PFkLfs1QcvL2gCKe6ElAGBP6TmIxgCQl0JDyavyUkM+iREquGnlJqYzQyLGU7rpA1qo6Yz7KvBpj
xGfWhHo0QXKmqUAIlY38w1QmwB6RVh63qY5i4rWhlG4rNj6gyvos6aSqOrH6Rp7jYkCYTejq5ArD
USZRw8Xgk6zn4Hg3AeY7udcFdP6p9WnvlO8Ntid4cJc/bZib3u4dfl+UkQqPQkr8ItVycCqn8qLS
LryXtMavVYYNrYHmZ7QCx8sOch+tsrmdYNEx26i4s1lwh2UYGjX7cJKg9SiwVnDi85VkgrR97A50
VOodaJluYWmvJQ==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity FIFO_SC_HS_Top is
port(
  Data :  in std_logic_vector(7 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(7 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end FIFO_SC_HS_Top;
architecture beh of FIFO_SC_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~fifo_sc_hs.FIFO_SC_HS_Top\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(7 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(7 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.FIFO_SC_HS_Top\
port map(
  Clk => Clk,
  Reset => Reset,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(7 downto 0) => Data(7 downto 0),
  Empty => Empty,
  Full => Full,
  Q(7 downto 0) => Q(7 downto 0));
end beh;
