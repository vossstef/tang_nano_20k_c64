library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.numeric_std.ALL;

package keyboard_matrix_pkg is
  type keyboard_t is array(14 downto 0, 7 downto 0) of std_logic;
end keyboard_matrix_pkg;  --end of package.

package body keyboard_matrix_pkg is

end keyboard_matrix_pkg; --end of the package body



