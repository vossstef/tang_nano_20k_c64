--
--Written by GowinSynthesis
--Product Version "V1.9.9 Beta-4 Education"
--Tue Apr 30 14:28:51 2024

--Source file index table:
--file0 "\/home/vossstef/Dokumente/gw_projects/tang_nano_20k_c64_dev/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\/home/vossstef/Dokumente/gw_projects/tang_nano_20k_c64_dev/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\/home/vossstef/Gowin_V1.9.9Beta-4_Education/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\/home/vossstef/Gowin_V1.9.9Beta-4_Education/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
Z9W/Q5MGSK7wnSPUDFFWQz8OFIcCI5cvY/8vdjkf4K7ZDZjNPJg6lcrVWm2L2lw9C83sNZ5R3Kp8
2llw1I8gljjMiGucgjIiOyzzSp2D6gAjsThfiy8AFnFvJxviEu9EIlEaVbUU4yF213RNzuChxeRI
QMKgIWW2UfqRJI32xbxoJ0U7PTOM/ZogNViAYF0j0QvVEEboLxL57BaFliZDntnBy0UPGy6Psvj8
Al4qiHHSlj1EnidE7h1HDMKQyVWWrAYI3dtDHAZjJNFA4RUeZThwwrQYkh+T6SsaoaDwn+iVqBg9
BO4XiYuk/xvTSkQgiwIHu1OtS6ZfD6mclK+oIg==

`protect encoding=(enctype="base64", line_length=76, bytes=13488)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
uraZTI5B4xdzGUP5m1gap1wTm0uPD+juDtFWd5nxgWAajtbJmjrK1IEzsznYkOiJ3X6qrT2LH6iS
n4N0JCJqhBf09pgwBvig30xjDwRQp4G2HHzUgF1sdeuT1VBEGtuPBDoxaJbdAkXC4GzZ2RxezYWZ
J0kB0OJMaD/mRLP++PN0Gm90rmnobwTgIPVcoJOWw409mTi/zsowWwDbwsziOaRJ/KaNCQoFcvxd
1GzB/iIk+TEN/NMnv4EKHu4OAu+2noRE4E1RQ5GjmFIRVYCdBJkJkW/F1ECKWsSbEDyTCx58ZHbr
AJ6oxBcphMWqZDkuEoTa9bKk1CTObCNsgCoOQ6HAPHB7pYW3k6xltxUfwPUqOVWd7PdYvGy+Tykx
LnzOkxrEU8iQ9dkm4oCb0KA7A1Mi/Xg39nFxADnrltMOt0j2yrtXdAKUnQplG8OSaZsdP6At8pIN
+baFk7CG6yO5dSXCrpnztz0L7dN/NY7AdIHqSK8FyC31WR1v6VaG/piW5kh5EjFOHwOGijmcToKr
vXbNWl4nnHYqY9npkO7OiXf4b3X7EzGEQJqd6vdbzRnelLr6rEWw6m1hV4vOL8sMKkjJ42DTyryZ
brflscgHBxN/tZRHeuM8roZmpV9M9NrhR6nBW7ZTmps2y8gsxO96VEJ7PgCpYWACSYi5N+BdfZb9
hQ1xHQPGngKjgVAIWqSjLx9eFJ5Rq/noBEQVLksLI/U1PsI8qrHNdZEeyMmUard/egtX9lwhKf0p
kutfxNQX9O2kTG6iakdPwM8rvWrS+5US2Kz3TM9Cmdfa1Z4xDg7JEal/qnKR3jKiPmR1naB4GoUX
7iU3AIS2CJS/ns5Xh8Ps3O7QOL67nzBDCCfxPkvU8FhEX/lsVREqZIdbda0zXMsLYSjcJ9pes9e2
BZJdE3eKjP6IwA+X3AM9QQhaYSdbbUl4pfmwxFQyYD7KpzyM3DKEkWIswDP8IQ1bmP97imMinWGb
bMdCU/wwDGrIEUnwCR41mBY62AnqSmvCT2JlVvTXxdHX7NtQJVCxWDHJN01ihYS5xVOtl7tadi/i
3qiFuJXclFkI7SQlD+WbOm8vT6sIOymmsCKBTwaYG3Z3NveTgRdX+rNVKe57Bl/NyRQaNlUqCtlt
g5vq1wEiytZDtvAcwEvRBx68FnMY9j/axtQ0lphzr2nS1Jb5EUTdfdvtktwIi/SFEz4PshNyo41n
fOuAtJn6AsdNQByBEVluAvMDX2BGasdXMIalBZBMVbVSfaczYF5VwgKz1qVqXQgmzbGYiuRX2MJC
uTkUmh8d8MpajZlqn2+xcxx29MgMsIt7QPLbnB+qJr5hGM3NSmumiDNPxEEqqQfemxItKZYIVuT1
rrWU5Fiw6zCQS/K6Y2e5LrqNzd6Q2gWD4SbKYJstJ0jWhEIS+zf2kETMlcSJIJDn0kc09tsUkZRB
dGdFVWuKB+RuMa5cpTcwDmLCaMRIr2niQILuPZSOz/oSPuJWOWQRkr4LzJpHHgYIkYAwlDHkcHht
fLI5MlaSE5yr62d1cdwO/bcdTSLUAVTBowUrzgy+rltpIz2hSqYETw0PRcTYLSfgszM9yzZL/fJh
S2pJQ5jGR1oc/OWJh+b2nivajCjFN6nfIImw4+5xxbfd/po2w3/Pe+cKCtY953bigzidKDAr1Z9Q
6Q/GBbRSfADa4SJ4tc8MdM5kFqcVI2qkqrMvr8zx9j1z1CjxE+8/kNUfkwUIDJewbbJk4gbrilAp
vZTCJAOV0ESPZ5CwOXyWmFywmuqniw0UnrjuVrwPfiJ6FCpWGBXmZUBpzydnaFzp/CTNebK5Egdj
M6CQyQuNi7++fSLty8PRFQ6HfcxYKPVlBHusBLmY7f3gRd/eu7VdLKW6p9cMoRaq7GMyZJyBA+W3
w0npS1729tH+OZvykpH/8gdzaM+GI6TwrTCSDlXXbowK1G2HtHpAaqaXkl5sBP/pM/yjS24ChTxe
v4yJbVtgeow+m8AQb6fwV5v9EglsI4Cl3FhyzsuRtlGI35vGjDWrNwc6b2vBwlNB4mNDoPtnafWQ
evaiSGRho8Rwx7wawQj4gH/TPiBtMu8YsBg6AxK4jYfVoha0rClQ0iEVsQghUdsBoNqIzNE3FlIR
qftU04lxUdeI2hnio62B1qy9o9WwHqc9VtqEhiNRuByJ8eEJggeWRY92FyCsMpBdCOdpKmo9lslb
rhppR93dbHVSdmbzBSWUi6dWdj9Y/Kv6GUdDCZH4LZauZ2tqmpjLAgL55jjSx/E5Kf9biufJAnd2
HTCp13zT39Bl+QhhpzAvD1Z9KyDGQbJjixZJLCQVcp1mGOJAANT3I+2Xs11sCqtKfsH3TgEdud/p
L4z5XlonufvhOJZ0p1Ap87M+ia9Ze0JYTXgiU11xNOhpnlbYtw7//YK1Udh/yBnpAWdUlbYvqHEI
qQU8B2HORfZhjIFJjzn20hRmLal0HxyyySGjt/zeEv03E46NRFlgBOFgF8zSb/CJL88P5RraQObS
rKKvOmZ7k7ccITXILOlP2WiFW7AG+w5+J5rDIrPZeEw2x+lBONBlivKQW3x1A9qj21yPEK76ID1w
8xiIJzR4SDUNHGgfZx3DsclXwD9Me+P+pPd4MOeC9D0qx1+4d2dn2nu4SeIC9t7Dvfq6tvvUlNoe
KslomBWSqDxvBkjwh1iYywcUb6pbTi2tnKUUVmgNDsLT31wf5h7+V++Z+el+Uv+/wwLCsj1RTTuw
s8kK1HonN0JbBiHxW9t2sOesNhUsEV+GMMQXrGlca5P0t/riAVEF/NLHiit3dvDULIrmE80M2OGt
Mzhw0czye2wjReuyxks3o2Owx7VdkbUaBG3GPmKwAwv54BUL+qgcXsFc/LJ9Ay1wPeEUtgqbR8LF
ST1E3CGYCX1zzSp+yArbEm8KthvWDoSKD3vzqXT0bZBTdNNBUPvl9fJ8KWCV0mhn7PGvwDv0FWgV
k347+rCnxWwaKcLZ+dnQ1QrdGtR5RrK1pmxbnVwQyZevMet1mJXG8/O5An/JHq1TPUiEqdH1qu1g
GLcvv4+uwpUGimdpwz/Eql4LPOPO805hXY0NEicsJTHzD5fyVhC7MI3UOwm5xb9Wi0c3ZBF93x3A
TDg9EprVoSQDDtiLiVex51ywstlXXGJapo6djmTYWumdDkK2TK2JzVyWQQAqN8bhgcUHr2A4JdxN
P//1TCGWrCaNJfSTdlYZcCL6H3yaHUX+5XEqtzf2z3VybtORo/pkbrAO7JcVvi+OQzFqXm71tTKT
XCSTsdtKYGKYJeHbqlk1IXSgAIyAteG4t7GQSIODOiJm+NQsFCZY+3qjCK+NGu1HARSqefr+XcKc
1ER5B5cxm8tN6QQ6hrw1dCYQBSBXBpW2bW1E+XkeutH5tH+3RSIeMGhiR+rvqstyBddclCxGL8iX
4M/4qZx7Fe9+3LlV2QI5Fe8vhx7VhCpyW1yOo6N/dwQnBMcaCR21dn8oTlHNqiT/ckohjzowJxWe
wRTsVvRj7z2cPdOu9ByIeLmYnk4/Ou5fUJ1sG+dJlr7WiTkNhY3itNnZKI28GeXj8MuupGAbrNU/
r//4kTb5ZrCHViAUwK16ibW3Kjdao1jTJM79v7VP3+j39jpoJo3/XbljYVxN8rp5eSf9GN5VstH1
7gUY4eNJyqkXQqdd50Fc+/vuaKuHF8Wsp18fSLewWwoZs4IB2jxXXeo8tzvBawrBlkMZTrtIDXVQ
H+i/qJ7+sd6cNyy5DbPvITZuuKcGamIf74V2iR0juwiAaJHrSJ7i/6peUbM/Y5HblwXe6jAe2V4K
a0SNEzSC6G0hyGOGn8OprmvRmITd7vDzxqemdD1EMlf8RHK06TJMOvQMSt/VLIh/wtqEIkgxQ5KJ
//W0lW6x6Pfaxo3H6tRzUuXbJGvm3sBgYkWwty8PdtV12eDjhhiPXcivQ0W/C2QrBj1nCk5pi3hk
VsTARFLUMEFQPg///1uoWJwCyj+GlH1t//5/PGU12GVhHWgSw0vSsLF5oSPgd9L/z/UZQDj3yM8Z
7VtRiKOpJiJBIbXB/nVGjZYEN3tsGNMazoCdR50UukMEuFeGaWrSBxtI3FAgUjoS38Zn6ZKk5cso
VTaZlCNvI898N5iCigyLfJdwZGxDziEpHBhG7GhTAhYyPUTCJEluW7nL2g/HUBgLliWq3HKrzjMo
qYIwVR0wxdCJJ+Rm+WTF7I31Tb/6v19O0zFlSH9YiZnt3+2NecHvHerTxBRdxGkEjb9GVzKRF95i
8M1JJfj+qP6bIC2MRGD2IdSnL1xy/FLQxCOvApiBJjnlUpzzpsxlo7Iodu/0mQTesmrflJakgN1o
DYOYWlVOOYlnt0Bducng5hS8C9qgPYMQT8bVizR285XTfJMJJmSPxGNjtN3NMgbAxK9iLqyCEYkI
hIEF7kLJQQrjbFpqb4wryaRep+ibBjxCJLqXwENfYniutsfvaYYtqbDClRAAvWvARBwPfbQmEFAz
1oJkN4yOO6GzuX7sau+w7/xKwef437mEMbOzKtXCDtRCZ5ivhPH99S2RZ2oZrg+OasYEdF/BwLVS
nUg4dbRrWZg4hzAzFI7GhvwMEhIgNXmjY6twBXgSKSMjBM1PC9N77wHpxktfyh0+UvVFT9liXoBl
7jv1lwPZhOsusM8DLiBzEHdwVRYIPArBAMu0tI+CiM3BeVACrg8zlnDR9LyBjYngLvlJHq5hXe5P
msNTEaJfDG+y3oRGNVPvFhpBHG9xeYlUDyRSo1ac3PzF0BXRH9QtEbM5FySgRBL9FRuBTV5Ow1Rt
StQWwDhxxHaoHVxesMt8JDv3dBdD/toaymKeudsyR8sSWhIt5CkrBe+Nf9cbHFPxPJJJ8fT4Z7Xa
5+IVDEyT6/czFsYvS+lxt8w9HwHBQK5+Rxi5Sxv3a76+U98QmveuUSr54h4UwkSpqPeCh6NLvs+/
vRU2NI8xY4vyO5WW0z5FXLj8HRMZGwEZg1QHjIqCQbJfnfrT/z4WboKPJNli8Av3LRsUVkwvBOWa
cfft+3rPUnTYOI4No1lglz50/MnHWh92j9S9dJy7ucMYXt1mtp3/+VTjAMa2doqdZOxTOJHAWuFZ
fJtehte1jKEL/g6D1UsL6yBUUNiJTqDQ6P16LFbxmOGcH+g7+uWa3fKI8s3fQX9kwSOv5QpTXa+x
XtB2lHjkzOvk+9dayQ1/OERWbIHRkOfxp/3b1j/Ve5xZl6EWEL0COheRekhFDkd8/evTm8qDNnI3
/cm8GsPPXWGLEUkFnJQuF3J5sxziwLhuKOW+8HUurqP9Z2DSBV+gIcY/ZG5xOjFLASHOaUvKgLsg
8cZcAZcIrm0QrsBTudtgiZoB94bV5SmjotM2uwY6EbGDYHYr1NM2XYDjZzmGrKEq1ExAwxh4VOH+
BukVkhJlLMQOoThKkRzIYaM6HTK8tOhcIPN4/0xf8advs5xyOsPooqWrnclkwXmZ+4gvXqpbE0nt
MW2Om83k3L0OH2RyJGEjDjV1/mA/MtzysysywrdSRRoWSS4eBbvzF6OLKAlsqAIChmSy0eV3SpUt
UNba5slXae9SzX3Amh/2N5VNbuO//+iM4LtnRyNuOZA5VmzshdatbURIvHwgDJ7GmtjVzECa0EMn
ddm//aV/IX8SBm0aahLSPx1t3ncNRInREZ8K9jIDv5dWPTwZtt7Yo462ARhi5daOTRcOQESL3Zc8
h2UrkkGf/RKc2vpzBPyCGsmjnrPbYcY0CRfC9A0bsJtpdBcJ+XFHJxkA31h0hrJQ33gO786Uc8lY
z5/01BUARgCqaStt3Pap1tWnTJV2H/vuuCXyHeeouBmjz0wZCQOMbousSpBpQO73sE/vfKbtCQmw
BDv1qJ1oQYMlovyhvAhxEaRRsxipoji9pJlX6OMK5sMeQLVoMtmF4EEMSV7vToDSG3rHjOLOHeI9
ZZbcbyDkTB87XFAJL+NN5FBNqy6dD+wJdna11E9JeOpqF8GhOwUviz5/FVEoNfdT77ToEtz8VXGO
LMgY0JlYmUodj6qGUhrgAN8RB6/wSVMTY9TJscyA606N/37qG3QkIzmsSibKPgezZdETrEXK4e/Q
mpKVGz1MHtDLaFbqGaVtRLPzvzcZHmm2f8bGMYNRHYjIfFFTDoTq73kejS3WiUzD/zpXYWtKQ1Lh
xVLMdNY/yvIYVpFw1A3T2ST369Fx+KORYxTWdFqo/bIs2Wv10yCFQHe0fuHQNSmtjwDXMCW3qksR
yNR+0knV5mEyaPHZhRK8GRcLnmtxkMmPjPzcTItxZM6xhS1/aohyHP3W2VHQewPV/DNxAZxpN6Qa
BWUUPE8CJ/45g27Mf5L99t77i5s64vVR3KmJOIRhgY+Nqf64FdPgEfKPDxyLLBofwZFMbkDItev0
33ic0kk9pWpafgXpc/M6X2ScemkANIvYJoFcKzFtHFFrWcEu7b7s7FNvFIZP5SbZRa4YpwwC+ePi
XFcyI11hBX/17DxFwng6h5P5LvAWvnPFkHcVff1KWgsqHxHeQmt4ORD+EPqz+2R7TtHnLDrW5PkK
l5uLvX21nXcXnNrkDZK6tObdd9FT2nVokQNZv5su4xXuYYCkB0ZUNYuIdEaQbE++L5Tcda86PFcW
m+2f7R1CcWFG5w0T2b2tZYAL00ueMF8YDYYWahXc2MFQZrTo5gWS63k93Coz13yDfcp0mdjTDSqz
dftNv0EF1A5cMeRYD0K9rk/GoQNT0PPfSeCaX0dSmGDvWgFCUBGMzQvCmBR8qiBt93YeJjvlqwkn
Fg1tjpmXJGpHtgtq/SsyYxwsOsIl3La5n42Fsud/yEsxsa+q9wmcM/XtqOYSGmlfse3P9OcV5ViL
60JvlLF5shq40DtxXfPQw3VtbLiUy3eraX3kwvApzjwrJE2OFshK3OWIBUqWWn/lRHQGtalS8cdj
Q8v8Q3JbkA12FVD/4mYwnjZNdbc5kW+axTTfzWWAQeHMSkXOID07UvgVFcSngdEGcuO31moKxnp7
KrPH4uo4KbiZTe8AqKvq/H6lkSHbytndDFtuoGbr+lD1EZrPKukNXxXxYP0Pw64e6NHpzawbjbuX
aUZJd38uGNMNM7i42hxbyOTvSZahuu9TAmF/TDkZAkCIeaph6AjmKOCZVNBRCUkOLG3rDMU8yx4V
mjiHxVPAi/P2ieyWmNYdizS0bnBg/J8MhdxWUck6eKIUWGX2LeUG4TqwQ47PzNSR3YVmzPZrIPzf
QifGPB6qbE73yzRYKl8mTEoEFpL8cEshSlegpS6CwgXfns5KU4JmVpF3cr+pESRB2mq+zRhJqZHJ
Si+TB9CqwTpWq4DAextPLO1vIMrDigk+0COCjiL7XGLk8jQ+8Pae0C+gykGy3zclJ6ZZ8oy45ZGx
vMFbf3pMb9WtAP4xqmDNfIHYyN7iCT1cKo3BPoQCpVywmG9EFdnsjezZHTWgq3KRnjwYTCgsxEab
9ZOAqRRjliZocX+a+/+Nn+KkiyWKPwWO5tCtaPi+l4icsruf/1AqVFal5d+DPgkNzkW5u3rEW0RR
pdoQXiU2FQ6wqdup2HUVTdJrxrmK/LFZuOPcVcE1WdDInu90nL9MY6QmaMFHR7IRUANgMs4kqgJl
gZ3/wG/IfTp8/ezsYh9VHIC4zGPpdGM5wYAwHQcUyr0lu34CHD6gvSeNaeZVM7oGfM4vxJa1hI9i
r7nokIydmP1W+RGovl2Qu1rEa0AnZOdIecBaybOA/RnxC0/O1wZZiT3rA73OLRwfDsgctHhux4tW
GMztmFdmElROlqKU0TrLTj/cT205M5MZgRQgaSRIyyK2k/ivdDCvLK2NcxFmMpdtcMvMU1b6tgZU
57s3p18Fvc2LQOOJDb2O6LaiL9AbZK2pz76bymEOqTbc584uUTU0wc9SREQZipdYjN6CHr2v6zW6
sVTazyFE7czzNO0JLta6ol9dKIujCQ+EHApRVcETOtB2n84HCsY8A/OePj9c+DHdGgXBNj8je6KE
zRd2kRea3t75kkYOV2RJWdHOBQWPGMquU1m8oqXzuMxg7o6Eu1833bVfPi1gkoWuLnSh+XGhN404
QKjVc6Ow3qDjr5Rgx/RkBx4oCXW3BDwURE9YQxMrexuDuWNe/kU+D+sbGB2M/5ho8qmGYVSpTNmf
F6s76iA3EkMNBPT5vf6mKU+sKQvafrwlXnbP7+lAkPD5qVyMw0Xq905o4HXxzaEAlGe7tyQLOSQv
ih//H0iyTAMQU3RdumitmKEQLF5MVKXnNmAG+pplEZI8HiGRQJwfhUFAbCuZGW8bFmxa7H7XepHs
OXmoWOcHjQG+mddzFLBm1c4HD0LrV1nRNQmCUdBqhpwLPS+lXcgiphrOsOmkOFM+Y79+PrnFfDD0
uIIbzyW0N2ZbPgZYLtahVy+y5JjIHFmxUq4qom6wI/qzl6+jRqstoG8cyoRAa3HruD8UyMwhBwY8
MAWEIRBBwL1oCh98lRxqem5XX2eRT/KpgrW51+SjG5ysb3BA9UVuxbuery6RVPD9nKJ8ndCFcKb2
trMZ7d7XvZLQ5zhMRE0y06g9rwhHM8T0BeK8RmpImaOc0xuPSCgjg3NTDSvSWI2PaCaMLpg40IFO
GwCfhkT9ucgaSXuv546SmZa9W8PSg52DZQoDJ4gfHATA0UUFw1t0/e70QlpANelZmZGWdMd7jTn3
ZTBR+BS9hwtt3IhJgeLyEeRDEjDJwAcX3lblZXkbfK6DBM31a3ZpbgopMo3aTw6Fp2duhF9ixbKR
i2OVyvqMYccC9nejAGp5sPJDp/BfbPRhHF6F0Zd3Izq9skudd3wj80YUjQTyagAEocR9jff/Ilir
I3XmZn/tULWcq3I6W4SqoLncCZw9Nm/bBkvnB6tZAqvjpEDh5GN1OQirpcrcI6X+vVLrYvhz3dmY
TyRv+0q32MAqSfkg1Rv/Rb7/xpsYISv7VK5IDu2cRZ61PsN15Jm0Ql7uqnq7W53fhC7cmyiBcmbw
PgOJbNHt/YMv+Md1Ek3rY1hRgX1xyG1bP619oIOcapTtt/nxe3MSpMFJDiTrarGzja5J+TfnRuRZ
V6ego67jeHTcE7L2Bm4O0fxzsPHMxcO9QF3pz/J6gwAzyoWLP1MbKZl4/UzknXnsDlUdJtEaE8zT
B3f9snBl0K466DsdrcfsC9sE5wujar3ZVY5AIDPToXpi0fa5ICyr5MuDPky2rh/Wj4kOqEBIGtaL
RufwS4UlHT4BmPc4sf/CeepWRCV3A7yElki9OVZ5CMuODDaViIiifPxP48bhKt4WjPMVOvoe3xy8
wDgkVObzrT+yt3kEghM/WZzDh5SWX0JMEq9hxcWWfnQZXMOV9UH4X184BwOpCcEs1eugKtEjiMyn
fE+3D+FN2VqMzVgqdqvk/EAqsniCAMxg0jbe+CTbc+q44H8PU75GgfwjVMHtPsHWlLE92M/T4BoH
sdKqC6BvbgTDErwGaBjVeWyhXmRzmGvnzIGQJ7NdAtk2ApnwuNMq4BvQ0Xj+CS8SGbQvkvuwDLD1
jBX+Jav+zhN1FWREtIJvG/VYOMnqyc7d7FrdhJS8FpX4pIPfKBneITMECPl2N5OqEDc2S4OqqbHw
bp1I5EHGFmTchEEO/lixc6+ZyKyae6Zwm/w9cmbS8rf6pWqS6Zw3JxpQidNY2OcV3xakAQMi+LTZ
baM1qy/7b8f+Ro3zSMSpkWhRbbsYUhv4tyAE/fDzhMvawbfnWrZQK7osy72prq5sMD2zW6ZOh8oV
+N8ELo3OdP7/qDRx7LecTrZYFd2SWfb/oX2tZam74oUU0ZdAvyyhx1BLgPqa3QH2wqjoqz9XK2h2
4L1ax0ZczgLgnyFbM8IyN00X3HSh4QYAxrKGz8HMiJ+EqXd1ldLxfissZP8G6DrmnKFeudhCgF4g
VXZfA2eeDggIZUmfel6UmzY1VRekAiLzFaS31JIZXWfhbcrAdbkp+VtYrLL52lgPa4Xa9pLZz6Az
zzl3XAjel+BfXivYofTpH6xzkEQ+WEdMGPUMNlNPKrfN1qP9JI1cwLpCZgLrL3M6ANylxFSaQ6su
rlkIuzq4YJJjwRiBW6zL3qxxJl36onOreSBx9+NMFamlg4p7uEnrRyJEA39OfuqUt9IYpmuSRaIW
RqG29cvwHCJE9d0JdoSyXWfUYPO3H0vV28eAeKVjgQ5AKmeRTxvEGUY3OKg+8ReG0LlvomijtkTi
6UtOntro2qeCsDytuZcD3NfOYu09gKFVLVeDP3PEpIOG5vrqrlFaTluCPnkgb3R0PD3mUQoO/5dd
TIHPWioZAb39b8A8CAPksKcBKNeI48IU2zfOOGZsBJ6hEsWMFbXfzD8f1f6V45JSs9tdlW4vouKS
uUBYbxbEtPfRUiKLpU/kAfcOKD3JaSXZ7o7EytNQTMWKULALIVLZfhw9nb+5/h7J86bE/zdB86Y3
XEvlN5azmnV8K8APaQwbQ0m/8I3KS6IYUa6EgYy55Fcmp0X1h5ML1T4Nt93kpIF3NaVM8lIzAgIm
XXgTxxqUb+OGR/Z+3DI4jZx5DWShl2ajGtTB5tCC/XEjEgoQP4JS0BzMiJ3lu64LS/llsNpJ3pCF
MI4aQExkrsLZi0v4WDuFeujrOLJ8at2wN6qW3p/NImQPcLIFXkHXQcA4ckfVhm+woFaS8rnlfaB+
ps/mkkkYm+zTZcPsGaee0UJz8vlXvgJDAsNNH0JXUhU9mI4lsoNGHRoTN9kvvjgoZBGbqybcS/4Y
ke4zJrfMy03f37UZHXQWMI+Qe4Oe/nkRWhVWSLnwekefB9HBNoLOm/ZKcPt+QDmKW3cPYsQc/ZVF
IVhpn5VRunmpUsxwitF8RtB/bsh0Y8V5XMv4gF5o5O+vko/q4qvcexR1EetXc5VXBSdZT5mLACb5
odC0Qbi9i30cHWPS44tXxdRu0JSkwY9VEREr73vZgC+qRDrEScIlmGfOLYeVFtjHq+oyFdH2ZVnA
8Mt8K8/aZY08u/5V7hyaYYKG0KyVIu6EQXMkzuNwylNaBgkWiVTJ2IvaZLTdon/8WzlLiuT/DgbW
iVLpxrE0SC7kXSGe07zFP6VWay5GEngUTxVf8UkBKJmUWtrkpDt05Vxxc8F6ZgKpxvkuD30NDfVz
T7SBmur/zmb/uoPuGwQt0Wf8wWu5WSW5PtGaDDC598QvNNR9HbZuUf29xaWSbmGxrItHy93+gCwT
w0AvD//YNVPsf1rIbgHAWlZ/M7QyCCtapgwpzjWWQ4qyCWZ/vzpmqKmHnRGVWrm3DA/8uxrHX9HD
NiuyyYxbkVzr9OdJIoM9aiv0E+MgSIYNsLqMMCeJXtN2biSvGbBXoOaHblGKCcufnDXH528Xmq2D
tVy1Jm3ubZT2ssSsSyOuDl59k1tZ9f3eMhU6f1NveazYofC/MOvutP9sPWnbBywkSje2VPKHUxAR
haNNhFJQWfuYWLmMAB/L2y+ieLrqPWj64976mwEEevaL0299JAkxHlLcwzSHYeUecY2HkYlt1mSU
jG4byH1M/YVHBdcqPXufx4kqHUCDI2eYyoscDh2shFUYI1BpsU57lNzyBJqZuhUWuh2nqcSqdUux
8hTK/sbGn9xWTfGkPuFusKIUHGO0oOlmv70DeS7+ETZtInpv/dvWR8qr3twO8v9kZnTmgCtyYtQq
+WDkGBojdGT2UdGN32vPF1dGSQO3VUyVjgYuAsWyjs4+4n7Cz7Iyz1FaHYrTl3WmML1i4Baqm6YU
8zsXEg3T1hvSBubOXYpUeDyJ7KQH0PagqwMHhY5zS/3rFtvZ2BQqvqWzewQqut1BnlGjL08pfyte
JMT4TyeV3xVefaSMgnSZTyQ4OxW3vntP6v+a5fekkDV7kPx5To2kOp9Dn5HJ2xkG2jfb3dT4lwIy
tQVCHYwFVqoNHzA5ZD7Kz8GQzLt7HqC9hio3WrcLnlO63x4fJCqFBBDmdyStmv5UWaYJ20RSz/78
lxD5CuhZc8y0j5obF7FVHz8doHepY7th/GTOX8TWNl7sr2FBeErd1ipt+G8xmXwn1oDSDNyP7RaO
6TOqwvHn3PmUrvRY9gvr3k9CbLrdaELczk8zsODcePz14PM8vijGJC0FYPKwiLvq+9IzTSC5LzeF
Ng0vdboh8XD3EjTCLmXxBM6crbV406Q909Ty20bpgGLQZiI17lWfKt2+mdh4mr9uxfk0o9ePrVVr
aG/GgsLqsuTcOku2uGwJj46PCEhQjdFbbk6Ny21910LyWAPUu2TzjNX/Z2RbQY7xa7lQ7s4d42EQ
iylDkiGgCVsGN7X4RL1MSVhIkHP5UADo0EqKx0pkVYWE57AzrD7VxiSE6yexgzBOQa8/QC/T1wFE
UpBs4BPgP4tlJ1MLFaNeJGnn1yj5rYaenhKX5Jlti3QIfnT8kD44UNG8gG8xdXayDfgHRGkKqm2s
3A3Iq6l8iddbRP0jnjRj538c7BY3jSuxNNgO+OJQ0E07aeabiU8cxmqoLh6JxgG0E9H444ZX4wfy
zuXG+PPsZ0OEoe1kABcXUcxw8SeRhZqCI1KmHtxBRlBrGSseKqLHXUyLtIKbknA4AFgEEtkqTL4y
owHWp6wQJtBDZhNQUnpKcpgZByrQGVmHcONP1CRcTqZxwI7FN+iwCj5Y0zjzDI3STVgKbFOts22a
0vq+/5GBkKjArxEwudyzHBWEYu95Z5aJFpPwsjHL/pJnLqO0AzZOl1njNZvNYG/yS07OZo2ZQgJw
GEbc9jHwakjOnn4qUAvyuJRLrHIxbX/luH4OWIpDLJ2NFnFi5Np/D2/SDKZsWnNTIXcTUhtbBcSl
kS6y3WZ7LOqhCggNsHA467lZqsLStcXLcL7DkjhP3hKTmdDYWdb+O8dYPqyDDe8PByrtexLJRHZO
Ubh9E1lkhPLgWul8z7fnhJbgLWQt5W/RLO57kR9NmO/EJRpFuxv23yMGlcPo6HCz76iDEK1h58nL
LnoPP93stEy2zDZFrDltZ0aG9ryyuIRaKKdAK1Dsq1KZ02ZKahLVxHmuuaRpdPhUF0rL041YKpxa
F6TalW8NsxQ5/4i+WGtFUVzrGQYoLAjw8Ie8IvZxuWILp5R1eZ1nAw5Y3slyK06aueS5jDrGhp8/
YjfZ2Zg3Z7f7OTXXk+RlWb1sZb0zjaSD2UOfzjKeHDVYTT+v6VVqdNaxgIvvgM5NKfT0gexSAD6H
/QPiBAn3zs/AP0JRbiPBKD1eVCZoKDRqISzm3QIQMGVMn7oj4Sf4sQTIQn/0qXPhSoxgihsPzEVE
fLSbuawy4iPVOKUQgjTbLTh9lbmc0gYUEleBjOhGKykB7THresjTNcP0CHf1B1oCPXp4sryh5ES6
OuaLT2I4+K2B5F8PhNuU/Ayx6lxjuTxUWMt0DL+RpFZ2GSjAg1fGJK1M0BKUuN4jgusTRVqH11IA
XQl4t5eqJxK4cjltCJvwZOH/N29KgvpR+ScgiP0XVvSnQdzBfD0q/5kNt2+7EC2RtuoztgK3yGde
GJpOYb2IbHCBpTw6EakTv4RoDKLUrKOpyqfxaMd59AJ92oj0lPy0D61IjDfSU6RXUPdFxXd8QJ9Y
yvof6c+NltJM+2Ft2UjrWAIvyixH2sPcjs8sEhZnC4jCQckk5ZGetrQewOMrDYOcGM/0d0cwyWRE
luJzzmQttG62eaL9Z8LGI1mh9VD/mNZARWNE/As9CWyxlFiHpIWQDjwm562864X9DRJaBhsbZ21w
veH5lZ23h3UvWvLlUaBBZf6Vw0PTHHgfwCyTfNS5cdJGo74D6wKhBX57Zd4hUEU8S8Qnbs+VCU8U
K/5tz2h5XYUx/8MUAMPUds+86pA00gyEP8QMJzmnittmW+FPmJgQAIxqwj5vU9fhiaLOxzTmoezM
CK9iYEHrfttJqwVJkMYP/K0U/e2Zt3OQ3zBlxtD6SzmqbmGyrR4Ag0+KKvTGF2OR+S0HB6/JRyIV
lPIr1MjAIpCmS53OA6hpcTAdLg6wa93a6yY4UAP4LOLpLq/rdQW+gQO02kHf9lAT2n2Xfi4gAXNG
J92RI8xmQSjizLbGyJK7SzkIJJBk1LZMrPh5v0Y5qkAjfIEKqc+YrYDkYQZ3MVUmifFDHpK4HQKQ
XmaizDPPFsl4gkgV/r5fQOhe6F/cVf78ZOLwK7ZtFmqsl5ONnaVsh0zcKitx+n5XdBkwNg0Vr1Hr
lvDW9lwto6DYUa4D5x/V7OIS/mzuktTjGS3fP48gGUAQEK0q/Hnz6+15PR5MntdkQT/Nqxa6dC+/
lTmSuHolcn7C0Ov83JSeIp4lvW3uN8k/F1hMcBkq64KlA4vqRY3bjd1n5pMXaekm9eSOzAMPwRal
FIzzGeB80jfNI0b/0ssNNY0Ca9q+T7O6UciLrMYi6y53sPkDLo/Q41iI6Uik+7ymU6ZatWtA5+3K
1E9iyR0Sj9N8RAcmrjt/TWQj4D8WzZSQQw13NIGhJvBzDIBxxbwZgmUDVb9ELobjakr9z/J0jqFL
2UkmVm5Vqlgn55rhGgzzPvnOOyG3EX5CiSv5yYCtNahh+4k5E68NTn6OhQzgF8KFeWDnwKYUIR+U
otuDGUWX4W7lo27ivezBYu4KUYqRgKiRViTq3uu1Wrzz5XpaObgYDwi3B3fgMUT5Ps7xFP9uK44q
j6pWrmUe5kFZY7ThunaFZRa5HFengxOm4bOrL0snpKvbsJffl7Wld+soVLqeZIJ696Nvsw5esguR
foPvGoI1Y7pK+ZBfSY05vMxBmZ/ootc27eFnAws9gMgg1xqAM/tv65pRJ1v1OfK7j5wO33UZleey
Q57LiIUlfsSgxm5E7ytPHcw/Tvq3QzhNRbvvgK1X84XiNGCuSECzR4iwpiiV6Qhz6s6ZiXraDm4E
0j5ROVDsW/w/3MZvxjSu4isdbZLOrTyYMXTokHJig+VYtrTt8c/JJXW8ASq1gNQzXr1gXTMcD6KV
4+2NJZWcHbzOBhqnp7BHwUsNkKpIxbTd3cMYFl5iXX7GawzEbQaFlPx9akBawmPf1ir+Ehlgq7Rl
Sf5bOAZi+Xj97FelwcCxc+RzZEHJ7BXAZ+b7jxAadJGmZxfQXwZSdqRag1p67zI7ICD1M+SFqkIg
fvFXC9WLtYM6kL6YmdvtcXoR3yMzUtICbLtFOG8V9SnT32x6CGcobZPXVVWCJqT/0MD1inicisWO
gzZw7WStXnkBxsuKHIG7udKnLaf052+rdyoDOO1Xz8HWyg8dy3RgiByZ4KomtC+eSqHeTl46zZYS
zsN2/iM+LtKsmgLOnFmz3swaNPyGcd37/6OGG5V+W7VqClN/iniWNK2zvXN6hHzmhRa4kzpHrPXt
kG9f0Heatf9rfDiwr6iaZ7umj9LMHadvPLY6E5vUeE1Ax1TVu4Lpj4E1XSsDDq8giPg2IfUYNbDd
xzzg8/3cXLxMr6JuOPzx57UYYdkTwom0CHyGHJHgRghcHKLDlznGCX8YSbuXnuBOXdyedTFgITOz
FODmkxkpCSiqFy/ZEIdIYY8njjTXiW8Fkj9YYsx8TjO6jneHl9Snd8HJWAAEfcPFSIUrcqSjixv6
+6maRZ26gQ5k7LaV+A3xQ0AXAJqBxbEoaeQozH+3Vuv4sNeA/qLM15sh9ytGF5ecPWNarYZati2c
1WA/9XTjoBKGFrXcTs6zgIbZKEnhDrCHjAPte4ZdwLOCklicUebowAlc7e4ZK/HQkBX3cmX8zMp8
/RfWHT2ICyB2VpyMPbw3NOcciAqqLTqzhSdUi6Ros95krY0alVbyTpoqxwve/ylc00zOvMq+2+fu
jv/DrtolGGivTK4oi16NXLXPDmYHP1zavhS8nAA1PYfbfQNoC7Vn4+Q33A+Xw9T7M8HYebZ7PNdl
nPaRyFqQiIZVybR7FghJrM90knGkdng2cq8cvwRHZ5pSb+uNxV/Dez0AjQX7ctxTAUCQjI3tbPHF
Tzzsh4EPpoecHHzTu5r8Hm/qlmaGSHaWyBx/y9StH4+unfMeqrPn5af/2tOGTHQLP5SSsBrL4g/Q
WMdWo8ifo60drGtnBhBn5Rzbj/PbkL33q5Dj9vq9sxY9T6twuU9FB10dh1VwrNo7+jEUpv/5+24b
vSmocIo6nL7zSf8n79OJgiswvjrE19jSbbZOXmgNf9GuDtmrwSyS89t3LxI5wVxnYThxHg8qRfoX
xSF3XOnMp9/83BcVLe68tBS5APJ0Nd0pmVwcnq4QFVWTNJ4NiErCEIDr6DacLFSY02JdvPaVsYPp
k4ODvLMrb88PX46BNrlXaDziXYS4lscr8B3j9DNSdtsLG9P9fuUi3KLVx+c+ijK5xf6FkslT34yg
uxSioPfaQOlhtfRPTRoispZTOkqloI7qia0Hi4ZQTwLbpwcy+lLa3m22esHCFhC3nZ3MPaJ1MK7q
fhmht8lS/Ci7v+Ii9WN9sKUoJgMbZhRmflWOCZuk3zkFWgB7dt6/k3AVcr/RzzRUHuaZ9mNfL0kp
0IOkFVxJU+AxZHCfd+r0bx9oZScPaVekWjTSrfSAfOSANxWRpCz55peLMgdMdAisUsytpuGzf1/1
ifz/YWtCCsz3R3NAeVpiqM8QpE7sG45cmTOxCmVbPwGTzaC801GYI5KjaJj+hxGzNxRe+h9d4TYB
4pPB9LGgzfGwKEXMqTs5CPRW3moSxkkKuW5YYHtROOc75UAQmUInmmQf05vnAGtlH/mmRjbrsxvG
1A7ws9ohla41EfgCllZIchmcSTKIJ5S0rbVJG0QMhfyO8lh8HKY/Xr0VbPfigIaFC2iGMJDbM9WJ
9OXysdDCC/HlKH5GOzEWNxJONTv8GgaYzh5wJUeErh+9rH+7LCe+ka5nMt7MfQMb856c8wQ82VKr
1B98FtjmpQun4kX4MFL4Se8XJheHH7IrG6l5TY1joXn9g++sEqjwCAvN61TugUsIymre2T8XoxXh
72daHWa9Q4Rr1Y8d7K9/axtaX4qwYhtWyqJhR41MNVMeVPLFKt5JQhWQJLw5jFQ70+mCl+iVUC0f
MMzfbs96rJoCNNGN0Gnb2EDRZvsEMddFgnNQaKKPib22jS+iuRDJYJVFtXXShkzw41xwdZmWI651
ghPKlhMQY0CHaHcXqIn9WQiVfsAlgmCK6hl7yZaJ+JhL8nImubYr/o/jNJoWH7KGj4yXTJXfGTzs
NLjQOJNtKP696GPblKq3K3TzGf+jIM/sbJqqBkayjzFuWg/OKUWsOnTm8W3Kq/4SU2B551vEgFin
9eGfrc4SAEDImtCZ/xPEDM+62upfbfqnVvBm3bkOjrV6IQN0pI0VT+Q64v1tA5/TAo1aH66LyojS
Zz+OiYQRnY4gIEhuBOAlZvpnBWvX3UlDoTby0bAp3aYO3GdYuB2OK5e+sFi/uAxnR6QLxh8nnTNN
FWCM5Fr376We1ZZ5iBkj4F9sbEPDJeldahy5ZLWGWRvdnmIvg0nNzEwW2ki5k7u1oFqMtua419o4
mwlt0Z9UMpBtrCtniVWQ10yV+9ucsqjw43wv9oshSULWCqBWVGNKnDlThAr57vvrgsSNiqWki5F6
sCFi9P0it/dHRTBpKDsX6EjWCRP1RGLyrbo29XWyajRsPB1Qsw4WgodoF905o19/lfJe3QoPDb0Q
8kYHpyuwHUrWN73n1ipYBAB+CGKoWRITupo34XtJLZVOhJrrXZKAjGZeokarVg+ma22GA00kjmhM
P9eUNe9hkaXcR26Wfy+4N/15VDBOuVmJSnkIIhgy+2Xvkaq9XYbQZkco5lwH9Yi5zbQ3dqKzCfv/
E9mbCSgj8dvXkeQ9xen3rlfA7qiL8NHyfy75D6L9hD6WZfDiixW6LdP5D5vAuSAl4gbXx9j7G11P
GnHQvWuBNlT1CuzvELibQxkQaI7VjwSz3ejqn6fVl0E8tlVyO+9+1qc/Wl3Av4pPoeat/4hm53I/
iAwl/QiSXaCOFDBsRrY2nvu7MEhgGcfAjLDR9DI8zk2wulOW3NRFV9BzJOCjbmzIgmEz0WXAORK5
Qy1qorSJoJROfY/bivchndpUaUuC+l/vqx0zdRXDkufY6JqC
`protect end_protected
