--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Thu Sep 07 20:15:52 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_RAM16S_color is
    port (
        dout: out std_logic_vector(3 downto 0);
        wre: in std_logic;
        ad: in std_logic_vector(9 downto 0);
        di: in std_logic_vector(3 downto 0);
        clk: in std_logic
    );
end Gowin_RAM16S_color;

architecture Behavioral of Gowin_RAM16S_color is

    signal ad4_inv: std_logic;
    signal ad5_inv: std_logic;
    signal ad6_inv: std_logic;
    signal lut_f_0: std_logic;
    signal ad7_inv: std_logic;
    signal ad8_inv: std_logic;
    signal ad9_inv: std_logic;
    signal lut_f_1: std_logic;
    signal lut_f_2: std_logic;
    signal lut_f_3: std_logic;
    signal lut_f_4: std_logic;
    signal lut_f_5: std_logic;
    signal lut_f_6: std_logic;
    signal lut_f_7: std_logic;
    signal lut_f_8: std_logic;
    signal lut_f_9: std_logic;
    signal lut_f_10: std_logic;
    signal lut_f_11: std_logic;
    signal lut_f_12: std_logic;
    signal lut_f_13: std_logic;
    signal lut_f_14: std_logic;
    signal lut_f_15: std_logic;
    signal lut_f_16: std_logic;
    signal lut_f_17: std_logic;
    signal lut_f_18: std_logic;
    signal lut_f_19: std_logic;
    signal lut_f_20: std_logic;
    signal lut_f_21: std_logic;
    signal lut_f_22: std_logic;
    signal lut_f_23: std_logic;
    signal lut_f_24: std_logic;
    signal lut_f_25: std_logic;
    signal lut_f_26: std_logic;
    signal lut_f_27: std_logic;
    signal lut_f_28: std_logic;
    signal lut_f_29: std_logic;
    signal lut_f_30: std_logic;
    signal lut_f_31: std_logic;
    signal lut_f_32: std_logic;
    signal lut_f_33: std_logic;
    signal lut_f_34: std_logic;
    signal lut_f_35: std_logic;
    signal lut_f_36: std_logic;
    signal lut_f_37: std_logic;
    signal lut_f_38: std_logic;
    signal lut_f_39: std_logic;
    signal lut_f_40: std_logic;
    signal lut_f_41: std_logic;
    signal lut_f_42: std_logic;
    signal lut_f_43: std_logic;
    signal lut_f_44: std_logic;
    signal lut_f_45: std_logic;
    signal lut_f_46: std_logic;
    signal lut_f_47: std_logic;
    signal lut_f_48: std_logic;
    signal lut_f_49: std_logic;
    signal lut_f_50: std_logic;
    signal lut_f_51: std_logic;
    signal lut_f_52: std_logic;
    signal lut_f_53: std_logic;
    signal lut_f_54: std_logic;
    signal lut_f_55: std_logic;
    signal lut_f_56: std_logic;
    signal lut_f_57: std_logic;
    signal lut_f_58: std_logic;
    signal lut_f_59: std_logic;
    signal lut_f_60: std_logic;
    signal lut_f_61: std_logic;
    signal lut_f_62: std_logic;
    signal lut_f_63: std_logic;
    signal lut_f_64: std_logic;
    signal lut_f_65: std_logic;
    signal lut_f_66: std_logic;
    signal lut_f_67: std_logic;
    signal lut_f_68: std_logic;
    signal lut_f_69: std_logic;
    signal lut_f_70: std_logic;
    signal lut_f_71: std_logic;
    signal lut_f_72: std_logic;
    signal lut_f_73: std_logic;
    signal lut_f_74: std_logic;
    signal lut_f_75: std_logic;
    signal lut_f_76: std_logic;
    signal lut_f_77: std_logic;
    signal lut_f_78: std_logic;
    signal lut_f_79: std_logic;
    signal lut_f_80: std_logic;
    signal lut_f_81: std_logic;
    signal lut_f_82: std_logic;
    signal lut_f_83: std_logic;
    signal lut_f_84: std_logic;
    signal lut_f_85: std_logic;
    signal lut_f_86: std_logic;
    signal lut_f_87: std_logic;
    signal lut_f_88: std_logic;
    signal lut_f_89: std_logic;
    signal lut_f_90: std_logic;
    signal lut_f_91: std_logic;
    signal lut_f_92: std_logic;
    signal lut_f_93: std_logic;
    signal lut_f_94: std_logic;
    signal lut_f_95: std_logic;
    signal lut_f_96: std_logic;
    signal lut_f_97: std_logic;
    signal lut_f_98: std_logic;
    signal lut_f_99: std_logic;
    signal lut_f_100: std_logic;
    signal lut_f_101: std_logic;
    signal lut_f_102: std_logic;
    signal lut_f_103: std_logic;
    signal lut_f_104: std_logic;
    signal lut_f_105: std_logic;
    signal lut_f_106: std_logic;
    signal lut_f_107: std_logic;
    signal lut_f_108: std_logic;
    signal lut_f_109: std_logic;
    signal lut_f_110: std_logic;
    signal lut_f_111: std_logic;
    signal lut_f_112: std_logic;
    signal lut_f_113: std_logic;
    signal lut_f_114: std_logic;
    signal lut_f_115: std_logic;
    signal lut_f_116: std_logic;
    signal lut_f_117: std_logic;
    signal lut_f_118: std_logic;
    signal lut_f_119: std_logic;
    signal lut_f_120: std_logic;
    signal lut_f_121: std_logic;
    signal lut_f_122: std_logic;
    signal lut_f_123: std_logic;
    signal lut_f_124: std_logic;
    signal lut_f_125: std_logic;
    signal lut_f_126: std_logic;
    signal lut_f_127: std_logic;
    signal ram16s_inst_0_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_1_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_2_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_3_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_4_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_5_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_6_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_7_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_8_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_9_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_10_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_11_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_12_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_13_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_14_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_15_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_16_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_17_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_18_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_19_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_20_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_21_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_22_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_23_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_24_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_25_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_26_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_27_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_28_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_29_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_30_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_31_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_32_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_33_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_34_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_35_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_36_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_37_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_38_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_39_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_40_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_41_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_42_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_43_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_44_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_45_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_46_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_47_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_48_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_49_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_50_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_51_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_52_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_53_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_54_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_55_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_56_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_57_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_58_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_59_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_60_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_61_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_62_dout: std_logic_vector(3 downto 0);
    signal ram16s_inst_63_dout: std_logic_vector(3 downto 0);
    signal mux_o_0: std_logic;
    signal mux_o_1: std_logic;
    signal mux_o_2: std_logic;
    signal mux_o_3: std_logic;
    signal mux_o_4: std_logic;
    signal mux_o_5: std_logic;
    signal mux_o_6: std_logic;
    signal mux_o_7: std_logic;
    signal mux_o_8: std_logic;
    signal mux_o_9: std_logic;
    signal mux_o_10: std_logic;
    signal mux_o_11: std_logic;
    signal mux_o_12: std_logic;
    signal mux_o_13: std_logic;
    signal mux_o_14: std_logic;
    signal mux_o_15: std_logic;
    signal mux_o_16: std_logic;
    signal mux_o_17: std_logic;
    signal mux_o_18: std_logic;
    signal mux_o_19: std_logic;
    signal mux_o_20: std_logic;
    signal mux_o_21: std_logic;
    signal mux_o_22: std_logic;
    signal mux_o_23: std_logic;
    signal mux_o_24: std_logic;
    signal mux_o_25: std_logic;
    signal mux_o_26: std_logic;
    signal mux_o_27: std_logic;
    signal mux_o_28: std_logic;
    signal mux_o_29: std_logic;
    signal mux_o_30: std_logic;
    signal mux_o_31: std_logic;
    signal mux_o_32: std_logic;
    signal mux_o_33: std_logic;
    signal mux_o_34: std_logic;
    signal mux_o_35: std_logic;
    signal mux_o_36: std_logic;
    signal mux_o_37: std_logic;
    signal mux_o_38: std_logic;
    signal mux_o_39: std_logic;
    signal mux_o_40: std_logic;
    signal mux_o_41: std_logic;
    signal mux_o_42: std_logic;
    signal mux_o_43: std_logic;
    signal mux_o_44: std_logic;
    signal mux_o_45: std_logic;
    signal mux_o_46: std_logic;
    signal mux_o_47: std_logic;
    signal mux_o_48: std_logic;
    signal mux_o_49: std_logic;
    signal mux_o_50: std_logic;
    signal mux_o_51: std_logic;
    signal mux_o_52: std_logic;
    signal mux_o_53: std_logic;
    signal mux_o_54: std_logic;
    signal mux_o_55: std_logic;
    signal mux_o_56: std_logic;
    signal mux_o_57: std_logic;
    signal mux_o_58: std_logic;
    signal mux_o_59: std_logic;
    signal mux_o_60: std_logic;
    signal mux_o_61: std_logic;
    signal mux_o_63: std_logic;
    signal mux_o_64: std_logic;
    signal mux_o_65: std_logic;
    signal mux_o_66: std_logic;
    signal mux_o_67: std_logic;
    signal mux_o_68: std_logic;
    signal mux_o_69: std_logic;
    signal mux_o_70: std_logic;
    signal mux_o_71: std_logic;
    signal mux_o_72: std_logic;
    signal mux_o_73: std_logic;
    signal mux_o_74: std_logic;
    signal mux_o_75: std_logic;
    signal mux_o_76: std_logic;
    signal mux_o_77: std_logic;
    signal mux_o_78: std_logic;
    signal mux_o_79: std_logic;
    signal mux_o_80: std_logic;
    signal mux_o_81: std_logic;
    signal mux_o_82: std_logic;
    signal mux_o_83: std_logic;
    signal mux_o_84: std_logic;
    signal mux_o_85: std_logic;
    signal mux_o_86: std_logic;
    signal mux_o_87: std_logic;
    signal mux_o_88: std_logic;
    signal mux_o_89: std_logic;
    signal mux_o_90: std_logic;
    signal mux_o_91: std_logic;
    signal mux_o_92: std_logic;
    signal mux_o_93: std_logic;
    signal mux_o_94: std_logic;
    signal mux_o_95: std_logic;
    signal mux_o_96: std_logic;
    signal mux_o_97: std_logic;
    signal mux_o_98: std_logic;
    signal mux_o_99: std_logic;
    signal mux_o_100: std_logic;
    signal mux_o_101: std_logic;
    signal mux_o_102: std_logic;
    signal mux_o_103: std_logic;
    signal mux_o_104: std_logic;
    signal mux_o_105: std_logic;
    signal mux_o_106: std_logic;
    signal mux_o_107: std_logic;
    signal mux_o_108: std_logic;
    signal mux_o_109: std_logic;
    signal mux_o_110: std_logic;
    signal mux_o_111: std_logic;
    signal mux_o_112: std_logic;
    signal mux_o_113: std_logic;
    signal mux_o_114: std_logic;
    signal mux_o_115: std_logic;
    signal mux_o_116: std_logic;
    signal mux_o_117: std_logic;
    signal mux_o_118: std_logic;
    signal mux_o_119: std_logic;
    signal mux_o_120: std_logic;
    signal mux_o_121: std_logic;
    signal mux_o_122: std_logic;
    signal mux_o_123: std_logic;
    signal mux_o_124: std_logic;
    signal mux_o_126: std_logic;
    signal mux_o_127: std_logic;
    signal mux_o_128: std_logic;
    signal mux_o_129: std_logic;
    signal mux_o_130: std_logic;
    signal mux_o_131: std_logic;
    signal mux_o_132: std_logic;
    signal mux_o_133: std_logic;
    signal mux_o_134: std_logic;
    signal mux_o_135: std_logic;
    signal mux_o_136: std_logic;
    signal mux_o_137: std_logic;
    signal mux_o_138: std_logic;
    signal mux_o_139: std_logic;
    signal mux_o_140: std_logic;
    signal mux_o_141: std_logic;
    signal mux_o_142: std_logic;
    signal mux_o_143: std_logic;
    signal mux_o_144: std_logic;
    signal mux_o_145: std_logic;
    signal mux_o_146: std_logic;
    signal mux_o_147: std_logic;
    signal mux_o_148: std_logic;
    signal mux_o_149: std_logic;
    signal mux_o_150: std_logic;
    signal mux_o_151: std_logic;
    signal mux_o_152: std_logic;
    signal mux_o_153: std_logic;
    signal mux_o_154: std_logic;
    signal mux_o_155: std_logic;
    signal mux_o_156: std_logic;
    signal mux_o_157: std_logic;
    signal mux_o_158: std_logic;
    signal mux_o_159: std_logic;
    signal mux_o_160: std_logic;
    signal mux_o_161: std_logic;
    signal mux_o_162: std_logic;
    signal mux_o_163: std_logic;
    signal mux_o_164: std_logic;
    signal mux_o_165: std_logic;
    signal mux_o_166: std_logic;
    signal mux_o_167: std_logic;
    signal mux_o_168: std_logic;
    signal mux_o_169: std_logic;
    signal mux_o_170: std_logic;
    signal mux_o_171: std_logic;
    signal mux_o_172: std_logic;
    signal mux_o_173: std_logic;
    signal mux_o_174: std_logic;
    signal mux_o_175: std_logic;
    signal mux_o_176: std_logic;
    signal mux_o_177: std_logic;
    signal mux_o_178: std_logic;
    signal mux_o_179: std_logic;
    signal mux_o_180: std_logic;
    signal mux_o_181: std_logic;
    signal mux_o_182: std_logic;
    signal mux_o_183: std_logic;
    signal mux_o_184: std_logic;
    signal mux_o_185: std_logic;
    signal mux_o_186: std_logic;
    signal mux_o_187: std_logic;
    signal mux_o_189: std_logic;
    signal mux_o_190: std_logic;
    signal mux_o_191: std_logic;
    signal mux_o_192: std_logic;
    signal mux_o_193: std_logic;
    signal mux_o_194: std_logic;
    signal mux_o_195: std_logic;
    signal mux_o_196: std_logic;
    signal mux_o_197: std_logic;
    signal mux_o_198: std_logic;
    signal mux_o_199: std_logic;
    signal mux_o_200: std_logic;
    signal mux_o_201: std_logic;
    signal mux_o_202: std_logic;
    signal mux_o_203: std_logic;
    signal mux_o_204: std_logic;
    signal mux_o_205: std_logic;
    signal mux_o_206: std_logic;
    signal mux_o_207: std_logic;
    signal mux_o_208: std_logic;
    signal mux_o_209: std_logic;
    signal mux_o_210: std_logic;
    signal mux_o_211: std_logic;
    signal mux_o_212: std_logic;
    signal mux_o_213: std_logic;
    signal mux_o_214: std_logic;
    signal mux_o_215: std_logic;
    signal mux_o_216: std_logic;
    signal mux_o_217: std_logic;
    signal mux_o_218: std_logic;
    signal mux_o_219: std_logic;
    signal mux_o_220: std_logic;
    signal mux_o_221: std_logic;
    signal mux_o_222: std_logic;
    signal mux_o_223: std_logic;
    signal mux_o_224: std_logic;
    signal mux_o_225: std_logic;
    signal mux_o_226: std_logic;
    signal mux_o_227: std_logic;
    signal mux_o_228: std_logic;
    signal mux_o_229: std_logic;
    signal mux_o_230: std_logic;
    signal mux_o_231: std_logic;
    signal mux_o_232: std_logic;
    signal mux_o_233: std_logic;
    signal mux_o_234: std_logic;
    signal mux_o_235: std_logic;
    signal mux_o_236: std_logic;
    signal mux_o_237: std_logic;
    signal mux_o_238: std_logic;
    signal mux_o_239: std_logic;
    signal mux_o_240: std_logic;
    signal mux_o_241: std_logic;
    signal mux_o_242: std_logic;
    signal mux_o_243: std_logic;
    signal mux_o_244: std_logic;
    signal mux_o_245: std_logic;
    signal mux_o_246: std_logic;
    signal mux_o_247: std_logic;
    signal mux_o_248: std_logic;
    signal mux_o_249: std_logic;
    signal mux_o_250: std_logic;

    -- component declaration
    component INV
        port (I: in std_logic; O: out std_logic);
    end component;

    -- component declaration
    component LUT4
        generic (
            INIT: in bit_vector := X"0000"
        );
        port (
            F: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            I2: in std_logic;
            I3: in std_logic
        );
    end component;

    --component declaration
    component RAM16S4
        GENERIC ( INIT_0 : bit_vector(15 downto 0) := X"0000";
                  INIT_1 : bit_vector(15 downto 0) := X"0000";
                  INIT_2 : bit_vector(15 downto 0) := X"0000";
                  INIT_3 : bit_vector(15 downto 0) := X"0000"
        );
        port (
            DO: out std_logic_vector(3 downto 0);
            DI: in std_logic_vector(3 downto 0);
            AD: in std_logic_vector(3 downto 0);
            WRE: in std_logic;
            CLK: in std_logic
        );
    end component;

    -- component declaration
    component MUX2
        port (
            O: out std_logic;
            I0: in std_logic;
            I1: in std_logic;
            S0: in std_logic
        );
    end component;

begin
    inv_inst_0 : INV
        port map (I => ad(4), O => ad4_inv);

    inv_inst_1 : INV
        port map (I => ad(5), O => ad5_inv);

    inv_inst_2 : INV
        port map (I => ad(6), O => ad6_inv);

    inv_inst_3 : INV
        port map (I => ad(7), O => ad7_inv);

    inv_inst_4 : INV
        port map (I => ad(8), O => ad8_inv);

    inv_inst_5 : INV
        port map (I => ad(9), O => ad9_inv);

    lut_inst_0 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_0,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_1 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_1,
            I0 => lut_f_0,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_2 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_2,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_3 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_3,
            I0 => lut_f_2,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_4 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_4,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_5 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_5,
            I0 => lut_f_4,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_6 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_6,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_7 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_7,
            I0 => lut_f_6,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_8 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_8,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_9 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_9,
            I0 => lut_f_8,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_10 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_10,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_11 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_11,
            I0 => lut_f_10,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_12 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_12,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_13 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_13,
            I0 => lut_f_12,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_14 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_14,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_15 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_15,
            I0 => lut_f_14,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_16 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_16,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_17 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_17,
            I0 => lut_f_16,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_18 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_18,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_19 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_19,
            I0 => lut_f_18,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_20 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_20,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_21 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_21,
            I0 => lut_f_20,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_22 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_22,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_23 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_23,
            I0 => lut_f_22,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_24 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_24,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_25 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_25,
            I0 => lut_f_24,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_26 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_26,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_27 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_27,
            I0 => lut_f_26,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_28 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_28,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_29 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_29,
            I0 => lut_f_28,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_30 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_30,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_31 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_31,
            I0 => lut_f_30,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad9_inv
        );

    lut_inst_32 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_32,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_33 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_33,
            I0 => lut_f_32,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_34 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_34,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_35 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_35,
            I0 => lut_f_34,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_36 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_36,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_37 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_37,
            I0 => lut_f_36,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_38 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_38,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_39 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_39,
            I0 => lut_f_38,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_40 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_40,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_41 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_41,
            I0 => lut_f_40,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_42 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_42,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_43 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_43,
            I0 => lut_f_42,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_44 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_44,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_45 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_45,
            I0 => lut_f_44,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_46 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_46,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_47 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_47,
            I0 => lut_f_46,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_48 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_48,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_49 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_49,
            I0 => lut_f_48,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_50 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_50,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_51 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_51,
            I0 => lut_f_50,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_52 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_52,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_53 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_53,
            I0 => lut_f_52,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_54 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_54,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_55 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_55,
            I0 => lut_f_54,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_56 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_56,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_57 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_57,
            I0 => lut_f_56,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_58 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_58,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_59 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_59,
            I0 => lut_f_58,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_60 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_60,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_61 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_61,
            I0 => lut_f_60,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_62 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_62,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_63 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_63,
            I0 => lut_f_62,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad9_inv
        );

    lut_inst_64 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_64,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_65 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_65,
            I0 => lut_f_64,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_66 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_66,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_67 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_67,
            I0 => lut_f_66,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_68 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_68,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_69 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_69,
            I0 => lut_f_68,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_70 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_70,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_71 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_71,
            I0 => lut_f_70,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_72 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_72,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_73 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_73,
            I0 => lut_f_72,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_74 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_74,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_75 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_75,
            I0 => lut_f_74,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_76 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_76,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_77 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_77,
            I0 => lut_f_76,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_78 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_78,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_79 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_79,
            I0 => lut_f_78,
            I1 => ad7_inv,
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_80 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_80,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_81 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_81,
            I0 => lut_f_80,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_82 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_82,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_83 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_83,
            I0 => lut_f_82,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_84 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_84,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_85 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_85,
            I0 => lut_f_84,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_86 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_86,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_87 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_87,
            I0 => lut_f_86,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_88 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_88,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_89 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_89,
            I0 => lut_f_88,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_90 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_90,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_91 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_91,
            I0 => lut_f_90,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_92 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_92,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_93 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_93,
            I0 => lut_f_92,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_94 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_94,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_95 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_95,
            I0 => lut_f_94,
            I1 => ad(7),
            I2 => ad8_inv,
            I3 => ad(9)
        );

    lut_inst_96 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_96,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_97 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_97,
            I0 => lut_f_96,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_98 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_98,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_99 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_99,
            I0 => lut_f_98,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_100 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_100,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_101 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_101,
            I0 => lut_f_100,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_102 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_102,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_103 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_103,
            I0 => lut_f_102,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_104 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_104,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_105 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_105,
            I0 => lut_f_104,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_106 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_106,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_107 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_107,
            I0 => lut_f_106,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_108 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_108,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_109 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_109,
            I0 => lut_f_108,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_110 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_110,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_111 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_111,
            I0 => lut_f_110,
            I1 => ad7_inv,
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_112 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_112,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_113 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_113,
            I0 => lut_f_112,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_114 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_114,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad6_inv
        );

    lut_inst_115 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_115,
            I0 => lut_f_114,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_116 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_116,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_117 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_117,
            I0 => lut_f_116,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_118 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_118,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad6_inv
        );

    lut_inst_119 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_119,
            I0 => lut_f_118,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_120 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_120,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_121 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_121,
            I0 => lut_f_120,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_122 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_122,
            I0 => wre,
            I1 => ad(4),
            I2 => ad5_inv,
            I3 => ad(6)
        );

    lut_inst_123 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_123,
            I0 => lut_f_122,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_124 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_124,
            I0 => wre,
            I1 => ad4_inv,
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_125 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_125,
            I0 => lut_f_124,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    lut_inst_126 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_126,
            I0 => wre,
            I1 => ad(4),
            I2 => ad(5),
            I3 => ad(6)
        );

    lut_inst_127 : LUT4
        generic map (
            INIT => X"8000"
        )
        port map (
            F => lut_f_127,
            I0 => lut_f_126,
            I1 => ad(7),
            I2 => ad(8),
            I3 => ad(9)
        );

    ram16s_inst_0: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_0_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_1,
            CLK => clk
        );

    ram16s_inst_1: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_1_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_3,
            CLK => clk
        );

    ram16s_inst_2: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_2_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_5,
            CLK => clk
        );

    ram16s_inst_3: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_3_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_7,
            CLK => clk
        );

    ram16s_inst_4: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_4_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_9,
            CLK => clk
        );

    ram16s_inst_5: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_5_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_11,
            CLK => clk
        );

    ram16s_inst_6: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_6_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_13,
            CLK => clk
        );

    ram16s_inst_7: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_7_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_15,
            CLK => clk
        );

    ram16s_inst_8: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_8_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_17,
            CLK => clk
        );

    ram16s_inst_9: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_9_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_19,
            CLK => clk
        );

    ram16s_inst_10: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_10_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_21,
            CLK => clk
        );

    ram16s_inst_11: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_11_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_23,
            CLK => clk
        );

    ram16s_inst_12: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_12_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_25,
            CLK => clk
        );

    ram16s_inst_13: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_13_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_27,
            CLK => clk
        );

    ram16s_inst_14: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_14_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_29,
            CLK => clk
        );

    ram16s_inst_15: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_15_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_31,
            CLK => clk
        );

    ram16s_inst_16: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_16_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_33,
            CLK => clk
        );

    ram16s_inst_17: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_17_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_35,
            CLK => clk
        );

    ram16s_inst_18: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_18_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_37,
            CLK => clk
        );

    ram16s_inst_19: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_19_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_39,
            CLK => clk
        );

    ram16s_inst_20: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_20_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_41,
            CLK => clk
        );

    ram16s_inst_21: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_21_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_43,
            CLK => clk
        );

    ram16s_inst_22: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_22_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_45,
            CLK => clk
        );

    ram16s_inst_23: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_23_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_47,
            CLK => clk
        );

    ram16s_inst_24: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_24_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_49,
            CLK => clk
        );

    ram16s_inst_25: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_25_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_51,
            CLK => clk
        );

    ram16s_inst_26: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_26_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_53,
            CLK => clk
        );

    ram16s_inst_27: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_27_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_55,
            CLK => clk
        );

    ram16s_inst_28: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_28_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_57,
            CLK => clk
        );

    ram16s_inst_29: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_29_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_59,
            CLK => clk
        );

    ram16s_inst_30: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_30_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_61,
            CLK => clk
        );

    ram16s_inst_31: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_31_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_63,
            CLK => clk
        );

    ram16s_inst_32: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_32_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_65,
            CLK => clk
        );

    ram16s_inst_33: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_33_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_67,
            CLK => clk
        );

    ram16s_inst_34: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_34_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_69,
            CLK => clk
        );

    ram16s_inst_35: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_35_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_71,
            CLK => clk
        );

    ram16s_inst_36: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_36_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_73,
            CLK => clk
        );

    ram16s_inst_37: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_37_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_75,
            CLK => clk
        );

    ram16s_inst_38: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_38_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_77,
            CLK => clk
        );

    ram16s_inst_39: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_39_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_79,
            CLK => clk
        );

    ram16s_inst_40: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_40_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_81,
            CLK => clk
        );

    ram16s_inst_41: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_41_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_83,
            CLK => clk
        );

    ram16s_inst_42: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_42_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_85,
            CLK => clk
        );

    ram16s_inst_43: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_43_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_87,
            CLK => clk
        );

    ram16s_inst_44: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_44_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_89,
            CLK => clk
        );

    ram16s_inst_45: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_45_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_91,
            CLK => clk
        );

    ram16s_inst_46: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_46_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_93,
            CLK => clk
        );

    ram16s_inst_47: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_47_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_95,
            CLK => clk
        );

    ram16s_inst_48: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_48_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_97,
            CLK => clk
        );

    ram16s_inst_49: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_49_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_99,
            CLK => clk
        );

    ram16s_inst_50: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_50_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_101,
            CLK => clk
        );

    ram16s_inst_51: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_51_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_103,
            CLK => clk
        );

    ram16s_inst_52: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_52_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_105,
            CLK => clk
        );

    ram16s_inst_53: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_53_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_107,
            CLK => clk
        );

    ram16s_inst_54: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_54_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_109,
            CLK => clk
        );

    ram16s_inst_55: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_55_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_111,
            CLK => clk
        );

    ram16s_inst_56: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_56_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_113,
            CLK => clk
        );

    ram16s_inst_57: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_57_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_115,
            CLK => clk
        );

    ram16s_inst_58: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_58_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_117,
            CLK => clk
        );

    ram16s_inst_59: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_59_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_119,
            CLK => clk
        );

    ram16s_inst_60: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_60_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_121,
            CLK => clk
        );

    ram16s_inst_61: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_61_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_123,
            CLK => clk
        );

    ram16s_inst_62: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_62_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_125,
            CLK => clk
        );

    ram16s_inst_63: RAM16S4
        generic map (
            INIT_0 => X"0000",
            INIT_1 => X"0000",
            INIT_2 => X"0000",
            INIT_3 => X"0000"
        )
        port map (
            DO => ram16s_inst_63_dout(3 downto 0),
            DI => di(3 downto 0),
            AD => ad(3 downto 0),
            WRE => lut_f_127,
            CLK => clk
        );

    mux_inst_0: MUX2
        port map (
            O => mux_o_0,
            I0 => ram16s_inst_0_dout(0),
            I1 => ram16s_inst_1_dout(0),
            S0 => ad(4)
        );

    mux_inst_1: MUX2
        port map (
            O => mux_o_1,
            I0 => ram16s_inst_2_dout(0),
            I1 => ram16s_inst_3_dout(0),
            S0 => ad(4)
        );

    mux_inst_2: MUX2
        port map (
            O => mux_o_2,
            I0 => ram16s_inst_4_dout(0),
            I1 => ram16s_inst_5_dout(0),
            S0 => ad(4)
        );

    mux_inst_3: MUX2
        port map (
            O => mux_o_3,
            I0 => ram16s_inst_6_dout(0),
            I1 => ram16s_inst_7_dout(0),
            S0 => ad(4)
        );

    mux_inst_4: MUX2
        port map (
            O => mux_o_4,
            I0 => ram16s_inst_8_dout(0),
            I1 => ram16s_inst_9_dout(0),
            S0 => ad(4)
        );

    mux_inst_5: MUX2
        port map (
            O => mux_o_5,
            I0 => ram16s_inst_10_dout(0),
            I1 => ram16s_inst_11_dout(0),
            S0 => ad(4)
        );

    mux_inst_6: MUX2
        port map (
            O => mux_o_6,
            I0 => ram16s_inst_12_dout(0),
            I1 => ram16s_inst_13_dout(0),
            S0 => ad(4)
        );

    mux_inst_7: MUX2
        port map (
            O => mux_o_7,
            I0 => ram16s_inst_14_dout(0),
            I1 => ram16s_inst_15_dout(0),
            S0 => ad(4)
        );

    mux_inst_8: MUX2
        port map (
            O => mux_o_8,
            I0 => ram16s_inst_16_dout(0),
            I1 => ram16s_inst_17_dout(0),
            S0 => ad(4)
        );

    mux_inst_9: MUX2
        port map (
            O => mux_o_9,
            I0 => ram16s_inst_18_dout(0),
            I1 => ram16s_inst_19_dout(0),
            S0 => ad(4)
        );

    mux_inst_10: MUX2
        port map (
            O => mux_o_10,
            I0 => ram16s_inst_20_dout(0),
            I1 => ram16s_inst_21_dout(0),
            S0 => ad(4)
        );

    mux_inst_11: MUX2
        port map (
            O => mux_o_11,
            I0 => ram16s_inst_22_dout(0),
            I1 => ram16s_inst_23_dout(0),
            S0 => ad(4)
        );

    mux_inst_12: MUX2
        port map (
            O => mux_o_12,
            I0 => ram16s_inst_24_dout(0),
            I1 => ram16s_inst_25_dout(0),
            S0 => ad(4)
        );

    mux_inst_13: MUX2
        port map (
            O => mux_o_13,
            I0 => ram16s_inst_26_dout(0),
            I1 => ram16s_inst_27_dout(0),
            S0 => ad(4)
        );

    mux_inst_14: MUX2
        port map (
            O => mux_o_14,
            I0 => ram16s_inst_28_dout(0),
            I1 => ram16s_inst_29_dout(0),
            S0 => ad(4)
        );

    mux_inst_15: MUX2
        port map (
            O => mux_o_15,
            I0 => ram16s_inst_30_dout(0),
            I1 => ram16s_inst_31_dout(0),
            S0 => ad(4)
        );

    mux_inst_16: MUX2
        port map (
            O => mux_o_16,
            I0 => ram16s_inst_32_dout(0),
            I1 => ram16s_inst_33_dout(0),
            S0 => ad(4)
        );

    mux_inst_17: MUX2
        port map (
            O => mux_o_17,
            I0 => ram16s_inst_34_dout(0),
            I1 => ram16s_inst_35_dout(0),
            S0 => ad(4)
        );

    mux_inst_18: MUX2
        port map (
            O => mux_o_18,
            I0 => ram16s_inst_36_dout(0),
            I1 => ram16s_inst_37_dout(0),
            S0 => ad(4)
        );

    mux_inst_19: MUX2
        port map (
            O => mux_o_19,
            I0 => ram16s_inst_38_dout(0),
            I1 => ram16s_inst_39_dout(0),
            S0 => ad(4)
        );

    mux_inst_20: MUX2
        port map (
            O => mux_o_20,
            I0 => ram16s_inst_40_dout(0),
            I1 => ram16s_inst_41_dout(0),
            S0 => ad(4)
        );

    mux_inst_21: MUX2
        port map (
            O => mux_o_21,
            I0 => ram16s_inst_42_dout(0),
            I1 => ram16s_inst_43_dout(0),
            S0 => ad(4)
        );

    mux_inst_22: MUX2
        port map (
            O => mux_o_22,
            I0 => ram16s_inst_44_dout(0),
            I1 => ram16s_inst_45_dout(0),
            S0 => ad(4)
        );

    mux_inst_23: MUX2
        port map (
            O => mux_o_23,
            I0 => ram16s_inst_46_dout(0),
            I1 => ram16s_inst_47_dout(0),
            S0 => ad(4)
        );

    mux_inst_24: MUX2
        port map (
            O => mux_o_24,
            I0 => ram16s_inst_48_dout(0),
            I1 => ram16s_inst_49_dout(0),
            S0 => ad(4)
        );

    mux_inst_25: MUX2
        port map (
            O => mux_o_25,
            I0 => ram16s_inst_50_dout(0),
            I1 => ram16s_inst_51_dout(0),
            S0 => ad(4)
        );

    mux_inst_26: MUX2
        port map (
            O => mux_o_26,
            I0 => ram16s_inst_52_dout(0),
            I1 => ram16s_inst_53_dout(0),
            S0 => ad(4)
        );

    mux_inst_27: MUX2
        port map (
            O => mux_o_27,
            I0 => ram16s_inst_54_dout(0),
            I1 => ram16s_inst_55_dout(0),
            S0 => ad(4)
        );

    mux_inst_28: MUX2
        port map (
            O => mux_o_28,
            I0 => ram16s_inst_56_dout(0),
            I1 => ram16s_inst_57_dout(0),
            S0 => ad(4)
        );

    mux_inst_29: MUX2
        port map (
            O => mux_o_29,
            I0 => ram16s_inst_58_dout(0),
            I1 => ram16s_inst_59_dout(0),
            S0 => ad(4)
        );

    mux_inst_30: MUX2
        port map (
            O => mux_o_30,
            I0 => ram16s_inst_60_dout(0),
            I1 => ram16s_inst_61_dout(0),
            S0 => ad(4)
        );

    mux_inst_31: MUX2
        port map (
            O => mux_o_31,
            I0 => ram16s_inst_62_dout(0),
            I1 => ram16s_inst_63_dout(0),
            S0 => ad(4)
        );

    mux_inst_32: MUX2
        port map (
            O => mux_o_32,
            I0 => mux_o_0,
            I1 => mux_o_1,
            S0 => ad(5)
        );

    mux_inst_33: MUX2
        port map (
            O => mux_o_33,
            I0 => mux_o_2,
            I1 => mux_o_3,
            S0 => ad(5)
        );

    mux_inst_34: MUX2
        port map (
            O => mux_o_34,
            I0 => mux_o_4,
            I1 => mux_o_5,
            S0 => ad(5)
        );

    mux_inst_35: MUX2
        port map (
            O => mux_o_35,
            I0 => mux_o_6,
            I1 => mux_o_7,
            S0 => ad(5)
        );

    mux_inst_36: MUX2
        port map (
            O => mux_o_36,
            I0 => mux_o_8,
            I1 => mux_o_9,
            S0 => ad(5)
        );

    mux_inst_37: MUX2
        port map (
            O => mux_o_37,
            I0 => mux_o_10,
            I1 => mux_o_11,
            S0 => ad(5)
        );

    mux_inst_38: MUX2
        port map (
            O => mux_o_38,
            I0 => mux_o_12,
            I1 => mux_o_13,
            S0 => ad(5)
        );

    mux_inst_39: MUX2
        port map (
            O => mux_o_39,
            I0 => mux_o_14,
            I1 => mux_o_15,
            S0 => ad(5)
        );

    mux_inst_40: MUX2
        port map (
            O => mux_o_40,
            I0 => mux_o_16,
            I1 => mux_o_17,
            S0 => ad(5)
        );

    mux_inst_41: MUX2
        port map (
            O => mux_o_41,
            I0 => mux_o_18,
            I1 => mux_o_19,
            S0 => ad(5)
        );

    mux_inst_42: MUX2
        port map (
            O => mux_o_42,
            I0 => mux_o_20,
            I1 => mux_o_21,
            S0 => ad(5)
        );

    mux_inst_43: MUX2
        port map (
            O => mux_o_43,
            I0 => mux_o_22,
            I1 => mux_o_23,
            S0 => ad(5)
        );

    mux_inst_44: MUX2
        port map (
            O => mux_o_44,
            I0 => mux_o_24,
            I1 => mux_o_25,
            S0 => ad(5)
        );

    mux_inst_45: MUX2
        port map (
            O => mux_o_45,
            I0 => mux_o_26,
            I1 => mux_o_27,
            S0 => ad(5)
        );

    mux_inst_46: MUX2
        port map (
            O => mux_o_46,
            I0 => mux_o_28,
            I1 => mux_o_29,
            S0 => ad(5)
        );

    mux_inst_47: MUX2
        port map (
            O => mux_o_47,
            I0 => mux_o_30,
            I1 => mux_o_31,
            S0 => ad(5)
        );

    mux_inst_48: MUX2
        port map (
            O => mux_o_48,
            I0 => mux_o_32,
            I1 => mux_o_33,
            S0 => ad(6)
        );

    mux_inst_49: MUX2
        port map (
            O => mux_o_49,
            I0 => mux_o_34,
            I1 => mux_o_35,
            S0 => ad(6)
        );

    mux_inst_50: MUX2
        port map (
            O => mux_o_50,
            I0 => mux_o_36,
            I1 => mux_o_37,
            S0 => ad(6)
        );

    mux_inst_51: MUX2
        port map (
            O => mux_o_51,
            I0 => mux_o_38,
            I1 => mux_o_39,
            S0 => ad(6)
        );

    mux_inst_52: MUX2
        port map (
            O => mux_o_52,
            I0 => mux_o_40,
            I1 => mux_o_41,
            S0 => ad(6)
        );

    mux_inst_53: MUX2
        port map (
            O => mux_o_53,
            I0 => mux_o_42,
            I1 => mux_o_43,
            S0 => ad(6)
        );

    mux_inst_54: MUX2
        port map (
            O => mux_o_54,
            I0 => mux_o_44,
            I1 => mux_o_45,
            S0 => ad(6)
        );

    mux_inst_55: MUX2
        port map (
            O => mux_o_55,
            I0 => mux_o_46,
            I1 => mux_o_47,
            S0 => ad(6)
        );

    mux_inst_56: MUX2
        port map (
            O => mux_o_56,
            I0 => mux_o_48,
            I1 => mux_o_49,
            S0 => ad(7)
        );

    mux_inst_57: MUX2
        port map (
            O => mux_o_57,
            I0 => mux_o_50,
            I1 => mux_o_51,
            S0 => ad(7)
        );

    mux_inst_58: MUX2
        port map (
            O => mux_o_58,
            I0 => mux_o_52,
            I1 => mux_o_53,
            S0 => ad(7)
        );

    mux_inst_59: MUX2
        port map (
            O => mux_o_59,
            I0 => mux_o_54,
            I1 => mux_o_55,
            S0 => ad(7)
        );

    mux_inst_60: MUX2
        port map (
            O => mux_o_60,
            I0 => mux_o_56,
            I1 => mux_o_57,
            S0 => ad(8)
        );

    mux_inst_61: MUX2
        port map (
            O => mux_o_61,
            I0 => mux_o_58,
            I1 => mux_o_59,
            S0 => ad(8)
        );

    mux_inst_62: MUX2
        port map (
            O => dout(0),
            I0 => mux_o_60,
            I1 => mux_o_61,
            S0 => ad(9)
        );

    mux_inst_63: MUX2
        port map (
            O => mux_o_63,
            I0 => ram16s_inst_0_dout(1),
            I1 => ram16s_inst_1_dout(1),
            S0 => ad(4)
        );

    mux_inst_64: MUX2
        port map (
            O => mux_o_64,
            I0 => ram16s_inst_2_dout(1),
            I1 => ram16s_inst_3_dout(1),
            S0 => ad(4)
        );

    mux_inst_65: MUX2
        port map (
            O => mux_o_65,
            I0 => ram16s_inst_4_dout(1),
            I1 => ram16s_inst_5_dout(1),
            S0 => ad(4)
        );

    mux_inst_66: MUX2
        port map (
            O => mux_o_66,
            I0 => ram16s_inst_6_dout(1),
            I1 => ram16s_inst_7_dout(1),
            S0 => ad(4)
        );

    mux_inst_67: MUX2
        port map (
            O => mux_o_67,
            I0 => ram16s_inst_8_dout(1),
            I1 => ram16s_inst_9_dout(1),
            S0 => ad(4)
        );

    mux_inst_68: MUX2
        port map (
            O => mux_o_68,
            I0 => ram16s_inst_10_dout(1),
            I1 => ram16s_inst_11_dout(1),
            S0 => ad(4)
        );

    mux_inst_69: MUX2
        port map (
            O => mux_o_69,
            I0 => ram16s_inst_12_dout(1),
            I1 => ram16s_inst_13_dout(1),
            S0 => ad(4)
        );

    mux_inst_70: MUX2
        port map (
            O => mux_o_70,
            I0 => ram16s_inst_14_dout(1),
            I1 => ram16s_inst_15_dout(1),
            S0 => ad(4)
        );

    mux_inst_71: MUX2
        port map (
            O => mux_o_71,
            I0 => ram16s_inst_16_dout(1),
            I1 => ram16s_inst_17_dout(1),
            S0 => ad(4)
        );

    mux_inst_72: MUX2
        port map (
            O => mux_o_72,
            I0 => ram16s_inst_18_dout(1),
            I1 => ram16s_inst_19_dout(1),
            S0 => ad(4)
        );

    mux_inst_73: MUX2
        port map (
            O => mux_o_73,
            I0 => ram16s_inst_20_dout(1),
            I1 => ram16s_inst_21_dout(1),
            S0 => ad(4)
        );

    mux_inst_74: MUX2
        port map (
            O => mux_o_74,
            I0 => ram16s_inst_22_dout(1),
            I1 => ram16s_inst_23_dout(1),
            S0 => ad(4)
        );

    mux_inst_75: MUX2
        port map (
            O => mux_o_75,
            I0 => ram16s_inst_24_dout(1),
            I1 => ram16s_inst_25_dout(1),
            S0 => ad(4)
        );

    mux_inst_76: MUX2
        port map (
            O => mux_o_76,
            I0 => ram16s_inst_26_dout(1),
            I1 => ram16s_inst_27_dout(1),
            S0 => ad(4)
        );

    mux_inst_77: MUX2
        port map (
            O => mux_o_77,
            I0 => ram16s_inst_28_dout(1),
            I1 => ram16s_inst_29_dout(1),
            S0 => ad(4)
        );

    mux_inst_78: MUX2
        port map (
            O => mux_o_78,
            I0 => ram16s_inst_30_dout(1),
            I1 => ram16s_inst_31_dout(1),
            S0 => ad(4)
        );

    mux_inst_79: MUX2
        port map (
            O => mux_o_79,
            I0 => ram16s_inst_32_dout(1),
            I1 => ram16s_inst_33_dout(1),
            S0 => ad(4)
        );

    mux_inst_80: MUX2
        port map (
            O => mux_o_80,
            I0 => ram16s_inst_34_dout(1),
            I1 => ram16s_inst_35_dout(1),
            S0 => ad(4)
        );

    mux_inst_81: MUX2
        port map (
            O => mux_o_81,
            I0 => ram16s_inst_36_dout(1),
            I1 => ram16s_inst_37_dout(1),
            S0 => ad(4)
        );

    mux_inst_82: MUX2
        port map (
            O => mux_o_82,
            I0 => ram16s_inst_38_dout(1),
            I1 => ram16s_inst_39_dout(1),
            S0 => ad(4)
        );

    mux_inst_83: MUX2
        port map (
            O => mux_o_83,
            I0 => ram16s_inst_40_dout(1),
            I1 => ram16s_inst_41_dout(1),
            S0 => ad(4)
        );

    mux_inst_84: MUX2
        port map (
            O => mux_o_84,
            I0 => ram16s_inst_42_dout(1),
            I1 => ram16s_inst_43_dout(1),
            S0 => ad(4)
        );

    mux_inst_85: MUX2
        port map (
            O => mux_o_85,
            I0 => ram16s_inst_44_dout(1),
            I1 => ram16s_inst_45_dout(1),
            S0 => ad(4)
        );

    mux_inst_86: MUX2
        port map (
            O => mux_o_86,
            I0 => ram16s_inst_46_dout(1),
            I1 => ram16s_inst_47_dout(1),
            S0 => ad(4)
        );

    mux_inst_87: MUX2
        port map (
            O => mux_o_87,
            I0 => ram16s_inst_48_dout(1),
            I1 => ram16s_inst_49_dout(1),
            S0 => ad(4)
        );

    mux_inst_88: MUX2
        port map (
            O => mux_o_88,
            I0 => ram16s_inst_50_dout(1),
            I1 => ram16s_inst_51_dout(1),
            S0 => ad(4)
        );

    mux_inst_89: MUX2
        port map (
            O => mux_o_89,
            I0 => ram16s_inst_52_dout(1),
            I1 => ram16s_inst_53_dout(1),
            S0 => ad(4)
        );

    mux_inst_90: MUX2
        port map (
            O => mux_o_90,
            I0 => ram16s_inst_54_dout(1),
            I1 => ram16s_inst_55_dout(1),
            S0 => ad(4)
        );

    mux_inst_91: MUX2
        port map (
            O => mux_o_91,
            I0 => ram16s_inst_56_dout(1),
            I1 => ram16s_inst_57_dout(1),
            S0 => ad(4)
        );

    mux_inst_92: MUX2
        port map (
            O => mux_o_92,
            I0 => ram16s_inst_58_dout(1),
            I1 => ram16s_inst_59_dout(1),
            S0 => ad(4)
        );

    mux_inst_93: MUX2
        port map (
            O => mux_o_93,
            I0 => ram16s_inst_60_dout(1),
            I1 => ram16s_inst_61_dout(1),
            S0 => ad(4)
        );

    mux_inst_94: MUX2
        port map (
            O => mux_o_94,
            I0 => ram16s_inst_62_dout(1),
            I1 => ram16s_inst_63_dout(1),
            S0 => ad(4)
        );

    mux_inst_95: MUX2
        port map (
            O => mux_o_95,
            I0 => mux_o_63,
            I1 => mux_o_64,
            S0 => ad(5)
        );

    mux_inst_96: MUX2
        port map (
            O => mux_o_96,
            I0 => mux_o_65,
            I1 => mux_o_66,
            S0 => ad(5)
        );

    mux_inst_97: MUX2
        port map (
            O => mux_o_97,
            I0 => mux_o_67,
            I1 => mux_o_68,
            S0 => ad(5)
        );

    mux_inst_98: MUX2
        port map (
            O => mux_o_98,
            I0 => mux_o_69,
            I1 => mux_o_70,
            S0 => ad(5)
        );

    mux_inst_99: MUX2
        port map (
            O => mux_o_99,
            I0 => mux_o_71,
            I1 => mux_o_72,
            S0 => ad(5)
        );

    mux_inst_100: MUX2
        port map (
            O => mux_o_100,
            I0 => mux_o_73,
            I1 => mux_o_74,
            S0 => ad(5)
        );

    mux_inst_101: MUX2
        port map (
            O => mux_o_101,
            I0 => mux_o_75,
            I1 => mux_o_76,
            S0 => ad(5)
        );

    mux_inst_102: MUX2
        port map (
            O => mux_o_102,
            I0 => mux_o_77,
            I1 => mux_o_78,
            S0 => ad(5)
        );

    mux_inst_103: MUX2
        port map (
            O => mux_o_103,
            I0 => mux_o_79,
            I1 => mux_o_80,
            S0 => ad(5)
        );

    mux_inst_104: MUX2
        port map (
            O => mux_o_104,
            I0 => mux_o_81,
            I1 => mux_o_82,
            S0 => ad(5)
        );

    mux_inst_105: MUX2
        port map (
            O => mux_o_105,
            I0 => mux_o_83,
            I1 => mux_o_84,
            S0 => ad(5)
        );

    mux_inst_106: MUX2
        port map (
            O => mux_o_106,
            I0 => mux_o_85,
            I1 => mux_o_86,
            S0 => ad(5)
        );

    mux_inst_107: MUX2
        port map (
            O => mux_o_107,
            I0 => mux_o_87,
            I1 => mux_o_88,
            S0 => ad(5)
        );

    mux_inst_108: MUX2
        port map (
            O => mux_o_108,
            I0 => mux_o_89,
            I1 => mux_o_90,
            S0 => ad(5)
        );

    mux_inst_109: MUX2
        port map (
            O => mux_o_109,
            I0 => mux_o_91,
            I1 => mux_o_92,
            S0 => ad(5)
        );

    mux_inst_110: MUX2
        port map (
            O => mux_o_110,
            I0 => mux_o_93,
            I1 => mux_o_94,
            S0 => ad(5)
        );

    mux_inst_111: MUX2
        port map (
            O => mux_o_111,
            I0 => mux_o_95,
            I1 => mux_o_96,
            S0 => ad(6)
        );

    mux_inst_112: MUX2
        port map (
            O => mux_o_112,
            I0 => mux_o_97,
            I1 => mux_o_98,
            S0 => ad(6)
        );

    mux_inst_113: MUX2
        port map (
            O => mux_o_113,
            I0 => mux_o_99,
            I1 => mux_o_100,
            S0 => ad(6)
        );

    mux_inst_114: MUX2
        port map (
            O => mux_o_114,
            I0 => mux_o_101,
            I1 => mux_o_102,
            S0 => ad(6)
        );

    mux_inst_115: MUX2
        port map (
            O => mux_o_115,
            I0 => mux_o_103,
            I1 => mux_o_104,
            S0 => ad(6)
        );

    mux_inst_116: MUX2
        port map (
            O => mux_o_116,
            I0 => mux_o_105,
            I1 => mux_o_106,
            S0 => ad(6)
        );

    mux_inst_117: MUX2
        port map (
            O => mux_o_117,
            I0 => mux_o_107,
            I1 => mux_o_108,
            S0 => ad(6)
        );

    mux_inst_118: MUX2
        port map (
            O => mux_o_118,
            I0 => mux_o_109,
            I1 => mux_o_110,
            S0 => ad(6)
        );

    mux_inst_119: MUX2
        port map (
            O => mux_o_119,
            I0 => mux_o_111,
            I1 => mux_o_112,
            S0 => ad(7)
        );

    mux_inst_120: MUX2
        port map (
            O => mux_o_120,
            I0 => mux_o_113,
            I1 => mux_o_114,
            S0 => ad(7)
        );

    mux_inst_121: MUX2
        port map (
            O => mux_o_121,
            I0 => mux_o_115,
            I1 => mux_o_116,
            S0 => ad(7)
        );

    mux_inst_122: MUX2
        port map (
            O => mux_o_122,
            I0 => mux_o_117,
            I1 => mux_o_118,
            S0 => ad(7)
        );

    mux_inst_123: MUX2
        port map (
            O => mux_o_123,
            I0 => mux_o_119,
            I1 => mux_o_120,
            S0 => ad(8)
        );

    mux_inst_124: MUX2
        port map (
            O => mux_o_124,
            I0 => mux_o_121,
            I1 => mux_o_122,
            S0 => ad(8)
        );

    mux_inst_125: MUX2
        port map (
            O => dout(1),
            I0 => mux_o_123,
            I1 => mux_o_124,
            S0 => ad(9)
        );

    mux_inst_126: MUX2
        port map (
            O => mux_o_126,
            I0 => ram16s_inst_0_dout(2),
            I1 => ram16s_inst_1_dout(2),
            S0 => ad(4)
        );

    mux_inst_127: MUX2
        port map (
            O => mux_o_127,
            I0 => ram16s_inst_2_dout(2),
            I1 => ram16s_inst_3_dout(2),
            S0 => ad(4)
        );

    mux_inst_128: MUX2
        port map (
            O => mux_o_128,
            I0 => ram16s_inst_4_dout(2),
            I1 => ram16s_inst_5_dout(2),
            S0 => ad(4)
        );

    mux_inst_129: MUX2
        port map (
            O => mux_o_129,
            I0 => ram16s_inst_6_dout(2),
            I1 => ram16s_inst_7_dout(2),
            S0 => ad(4)
        );

    mux_inst_130: MUX2
        port map (
            O => mux_o_130,
            I0 => ram16s_inst_8_dout(2),
            I1 => ram16s_inst_9_dout(2),
            S0 => ad(4)
        );

    mux_inst_131: MUX2
        port map (
            O => mux_o_131,
            I0 => ram16s_inst_10_dout(2),
            I1 => ram16s_inst_11_dout(2),
            S0 => ad(4)
        );

    mux_inst_132: MUX2
        port map (
            O => mux_o_132,
            I0 => ram16s_inst_12_dout(2),
            I1 => ram16s_inst_13_dout(2),
            S0 => ad(4)
        );

    mux_inst_133: MUX2
        port map (
            O => mux_o_133,
            I0 => ram16s_inst_14_dout(2),
            I1 => ram16s_inst_15_dout(2),
            S0 => ad(4)
        );

    mux_inst_134: MUX2
        port map (
            O => mux_o_134,
            I0 => ram16s_inst_16_dout(2),
            I1 => ram16s_inst_17_dout(2),
            S0 => ad(4)
        );

    mux_inst_135: MUX2
        port map (
            O => mux_o_135,
            I0 => ram16s_inst_18_dout(2),
            I1 => ram16s_inst_19_dout(2),
            S0 => ad(4)
        );

    mux_inst_136: MUX2
        port map (
            O => mux_o_136,
            I0 => ram16s_inst_20_dout(2),
            I1 => ram16s_inst_21_dout(2),
            S0 => ad(4)
        );

    mux_inst_137: MUX2
        port map (
            O => mux_o_137,
            I0 => ram16s_inst_22_dout(2),
            I1 => ram16s_inst_23_dout(2),
            S0 => ad(4)
        );

    mux_inst_138: MUX2
        port map (
            O => mux_o_138,
            I0 => ram16s_inst_24_dout(2),
            I1 => ram16s_inst_25_dout(2),
            S0 => ad(4)
        );

    mux_inst_139: MUX2
        port map (
            O => mux_o_139,
            I0 => ram16s_inst_26_dout(2),
            I1 => ram16s_inst_27_dout(2),
            S0 => ad(4)
        );

    mux_inst_140: MUX2
        port map (
            O => mux_o_140,
            I0 => ram16s_inst_28_dout(2),
            I1 => ram16s_inst_29_dout(2),
            S0 => ad(4)
        );

    mux_inst_141: MUX2
        port map (
            O => mux_o_141,
            I0 => ram16s_inst_30_dout(2),
            I1 => ram16s_inst_31_dout(2),
            S0 => ad(4)
        );

    mux_inst_142: MUX2
        port map (
            O => mux_o_142,
            I0 => ram16s_inst_32_dout(2),
            I1 => ram16s_inst_33_dout(2),
            S0 => ad(4)
        );

    mux_inst_143: MUX2
        port map (
            O => mux_o_143,
            I0 => ram16s_inst_34_dout(2),
            I1 => ram16s_inst_35_dout(2),
            S0 => ad(4)
        );

    mux_inst_144: MUX2
        port map (
            O => mux_o_144,
            I0 => ram16s_inst_36_dout(2),
            I1 => ram16s_inst_37_dout(2),
            S0 => ad(4)
        );

    mux_inst_145: MUX2
        port map (
            O => mux_o_145,
            I0 => ram16s_inst_38_dout(2),
            I1 => ram16s_inst_39_dout(2),
            S0 => ad(4)
        );

    mux_inst_146: MUX2
        port map (
            O => mux_o_146,
            I0 => ram16s_inst_40_dout(2),
            I1 => ram16s_inst_41_dout(2),
            S0 => ad(4)
        );

    mux_inst_147: MUX2
        port map (
            O => mux_o_147,
            I0 => ram16s_inst_42_dout(2),
            I1 => ram16s_inst_43_dout(2),
            S0 => ad(4)
        );

    mux_inst_148: MUX2
        port map (
            O => mux_o_148,
            I0 => ram16s_inst_44_dout(2),
            I1 => ram16s_inst_45_dout(2),
            S0 => ad(4)
        );

    mux_inst_149: MUX2
        port map (
            O => mux_o_149,
            I0 => ram16s_inst_46_dout(2),
            I1 => ram16s_inst_47_dout(2),
            S0 => ad(4)
        );

    mux_inst_150: MUX2
        port map (
            O => mux_o_150,
            I0 => ram16s_inst_48_dout(2),
            I1 => ram16s_inst_49_dout(2),
            S0 => ad(4)
        );

    mux_inst_151: MUX2
        port map (
            O => mux_o_151,
            I0 => ram16s_inst_50_dout(2),
            I1 => ram16s_inst_51_dout(2),
            S0 => ad(4)
        );

    mux_inst_152: MUX2
        port map (
            O => mux_o_152,
            I0 => ram16s_inst_52_dout(2),
            I1 => ram16s_inst_53_dout(2),
            S0 => ad(4)
        );

    mux_inst_153: MUX2
        port map (
            O => mux_o_153,
            I0 => ram16s_inst_54_dout(2),
            I1 => ram16s_inst_55_dout(2),
            S0 => ad(4)
        );

    mux_inst_154: MUX2
        port map (
            O => mux_o_154,
            I0 => ram16s_inst_56_dout(2),
            I1 => ram16s_inst_57_dout(2),
            S0 => ad(4)
        );

    mux_inst_155: MUX2
        port map (
            O => mux_o_155,
            I0 => ram16s_inst_58_dout(2),
            I1 => ram16s_inst_59_dout(2),
            S0 => ad(4)
        );

    mux_inst_156: MUX2
        port map (
            O => mux_o_156,
            I0 => ram16s_inst_60_dout(2),
            I1 => ram16s_inst_61_dout(2),
            S0 => ad(4)
        );

    mux_inst_157: MUX2
        port map (
            O => mux_o_157,
            I0 => ram16s_inst_62_dout(2),
            I1 => ram16s_inst_63_dout(2),
            S0 => ad(4)
        );

    mux_inst_158: MUX2
        port map (
            O => mux_o_158,
            I0 => mux_o_126,
            I1 => mux_o_127,
            S0 => ad(5)
        );

    mux_inst_159: MUX2
        port map (
            O => mux_o_159,
            I0 => mux_o_128,
            I1 => mux_o_129,
            S0 => ad(5)
        );

    mux_inst_160: MUX2
        port map (
            O => mux_o_160,
            I0 => mux_o_130,
            I1 => mux_o_131,
            S0 => ad(5)
        );

    mux_inst_161: MUX2
        port map (
            O => mux_o_161,
            I0 => mux_o_132,
            I1 => mux_o_133,
            S0 => ad(5)
        );

    mux_inst_162: MUX2
        port map (
            O => mux_o_162,
            I0 => mux_o_134,
            I1 => mux_o_135,
            S0 => ad(5)
        );

    mux_inst_163: MUX2
        port map (
            O => mux_o_163,
            I0 => mux_o_136,
            I1 => mux_o_137,
            S0 => ad(5)
        );

    mux_inst_164: MUX2
        port map (
            O => mux_o_164,
            I0 => mux_o_138,
            I1 => mux_o_139,
            S0 => ad(5)
        );

    mux_inst_165: MUX2
        port map (
            O => mux_o_165,
            I0 => mux_o_140,
            I1 => mux_o_141,
            S0 => ad(5)
        );

    mux_inst_166: MUX2
        port map (
            O => mux_o_166,
            I0 => mux_o_142,
            I1 => mux_o_143,
            S0 => ad(5)
        );

    mux_inst_167: MUX2
        port map (
            O => mux_o_167,
            I0 => mux_o_144,
            I1 => mux_o_145,
            S0 => ad(5)
        );

    mux_inst_168: MUX2
        port map (
            O => mux_o_168,
            I0 => mux_o_146,
            I1 => mux_o_147,
            S0 => ad(5)
        );

    mux_inst_169: MUX2
        port map (
            O => mux_o_169,
            I0 => mux_o_148,
            I1 => mux_o_149,
            S0 => ad(5)
        );

    mux_inst_170: MUX2
        port map (
            O => mux_o_170,
            I0 => mux_o_150,
            I1 => mux_o_151,
            S0 => ad(5)
        );

    mux_inst_171: MUX2
        port map (
            O => mux_o_171,
            I0 => mux_o_152,
            I1 => mux_o_153,
            S0 => ad(5)
        );

    mux_inst_172: MUX2
        port map (
            O => mux_o_172,
            I0 => mux_o_154,
            I1 => mux_o_155,
            S0 => ad(5)
        );

    mux_inst_173: MUX2
        port map (
            O => mux_o_173,
            I0 => mux_o_156,
            I1 => mux_o_157,
            S0 => ad(5)
        );

    mux_inst_174: MUX2
        port map (
            O => mux_o_174,
            I0 => mux_o_158,
            I1 => mux_o_159,
            S0 => ad(6)
        );

    mux_inst_175: MUX2
        port map (
            O => mux_o_175,
            I0 => mux_o_160,
            I1 => mux_o_161,
            S0 => ad(6)
        );

    mux_inst_176: MUX2
        port map (
            O => mux_o_176,
            I0 => mux_o_162,
            I1 => mux_o_163,
            S0 => ad(6)
        );

    mux_inst_177: MUX2
        port map (
            O => mux_o_177,
            I0 => mux_o_164,
            I1 => mux_o_165,
            S0 => ad(6)
        );

    mux_inst_178: MUX2
        port map (
            O => mux_o_178,
            I0 => mux_o_166,
            I1 => mux_o_167,
            S0 => ad(6)
        );

    mux_inst_179: MUX2
        port map (
            O => mux_o_179,
            I0 => mux_o_168,
            I1 => mux_o_169,
            S0 => ad(6)
        );

    mux_inst_180: MUX2
        port map (
            O => mux_o_180,
            I0 => mux_o_170,
            I1 => mux_o_171,
            S0 => ad(6)
        );

    mux_inst_181: MUX2
        port map (
            O => mux_o_181,
            I0 => mux_o_172,
            I1 => mux_o_173,
            S0 => ad(6)
        );

    mux_inst_182: MUX2
        port map (
            O => mux_o_182,
            I0 => mux_o_174,
            I1 => mux_o_175,
            S0 => ad(7)
        );

    mux_inst_183: MUX2
        port map (
            O => mux_o_183,
            I0 => mux_o_176,
            I1 => mux_o_177,
            S0 => ad(7)
        );

    mux_inst_184: MUX2
        port map (
            O => mux_o_184,
            I0 => mux_o_178,
            I1 => mux_o_179,
            S0 => ad(7)
        );

    mux_inst_185: MUX2
        port map (
            O => mux_o_185,
            I0 => mux_o_180,
            I1 => mux_o_181,
            S0 => ad(7)
        );

    mux_inst_186: MUX2
        port map (
            O => mux_o_186,
            I0 => mux_o_182,
            I1 => mux_o_183,
            S0 => ad(8)
        );

    mux_inst_187: MUX2
        port map (
            O => mux_o_187,
            I0 => mux_o_184,
            I1 => mux_o_185,
            S0 => ad(8)
        );

    mux_inst_188: MUX2
        port map (
            O => dout(2),
            I0 => mux_o_186,
            I1 => mux_o_187,
            S0 => ad(9)
        );

    mux_inst_189: MUX2
        port map (
            O => mux_o_189,
            I0 => ram16s_inst_0_dout(3),
            I1 => ram16s_inst_1_dout(3),
            S0 => ad(4)
        );

    mux_inst_190: MUX2
        port map (
            O => mux_o_190,
            I0 => ram16s_inst_2_dout(3),
            I1 => ram16s_inst_3_dout(3),
            S0 => ad(4)
        );

    mux_inst_191: MUX2
        port map (
            O => mux_o_191,
            I0 => ram16s_inst_4_dout(3),
            I1 => ram16s_inst_5_dout(3),
            S0 => ad(4)
        );

    mux_inst_192: MUX2
        port map (
            O => mux_o_192,
            I0 => ram16s_inst_6_dout(3),
            I1 => ram16s_inst_7_dout(3),
            S0 => ad(4)
        );

    mux_inst_193: MUX2
        port map (
            O => mux_o_193,
            I0 => ram16s_inst_8_dout(3),
            I1 => ram16s_inst_9_dout(3),
            S0 => ad(4)
        );

    mux_inst_194: MUX2
        port map (
            O => mux_o_194,
            I0 => ram16s_inst_10_dout(3),
            I1 => ram16s_inst_11_dout(3),
            S0 => ad(4)
        );

    mux_inst_195: MUX2
        port map (
            O => mux_o_195,
            I0 => ram16s_inst_12_dout(3),
            I1 => ram16s_inst_13_dout(3),
            S0 => ad(4)
        );

    mux_inst_196: MUX2
        port map (
            O => mux_o_196,
            I0 => ram16s_inst_14_dout(3),
            I1 => ram16s_inst_15_dout(3),
            S0 => ad(4)
        );

    mux_inst_197: MUX2
        port map (
            O => mux_o_197,
            I0 => ram16s_inst_16_dout(3),
            I1 => ram16s_inst_17_dout(3),
            S0 => ad(4)
        );

    mux_inst_198: MUX2
        port map (
            O => mux_o_198,
            I0 => ram16s_inst_18_dout(3),
            I1 => ram16s_inst_19_dout(3),
            S0 => ad(4)
        );

    mux_inst_199: MUX2
        port map (
            O => mux_o_199,
            I0 => ram16s_inst_20_dout(3),
            I1 => ram16s_inst_21_dout(3),
            S0 => ad(4)
        );

    mux_inst_200: MUX2
        port map (
            O => mux_o_200,
            I0 => ram16s_inst_22_dout(3),
            I1 => ram16s_inst_23_dout(3),
            S0 => ad(4)
        );

    mux_inst_201: MUX2
        port map (
            O => mux_o_201,
            I0 => ram16s_inst_24_dout(3),
            I1 => ram16s_inst_25_dout(3),
            S0 => ad(4)
        );

    mux_inst_202: MUX2
        port map (
            O => mux_o_202,
            I0 => ram16s_inst_26_dout(3),
            I1 => ram16s_inst_27_dout(3),
            S0 => ad(4)
        );

    mux_inst_203: MUX2
        port map (
            O => mux_o_203,
            I0 => ram16s_inst_28_dout(3),
            I1 => ram16s_inst_29_dout(3),
            S0 => ad(4)
        );

    mux_inst_204: MUX2
        port map (
            O => mux_o_204,
            I0 => ram16s_inst_30_dout(3),
            I1 => ram16s_inst_31_dout(3),
            S0 => ad(4)
        );

    mux_inst_205: MUX2
        port map (
            O => mux_o_205,
            I0 => ram16s_inst_32_dout(3),
            I1 => ram16s_inst_33_dout(3),
            S0 => ad(4)
        );

    mux_inst_206: MUX2
        port map (
            O => mux_o_206,
            I0 => ram16s_inst_34_dout(3),
            I1 => ram16s_inst_35_dout(3),
            S0 => ad(4)
        );

    mux_inst_207: MUX2
        port map (
            O => mux_o_207,
            I0 => ram16s_inst_36_dout(3),
            I1 => ram16s_inst_37_dout(3),
            S0 => ad(4)
        );

    mux_inst_208: MUX2
        port map (
            O => mux_o_208,
            I0 => ram16s_inst_38_dout(3),
            I1 => ram16s_inst_39_dout(3),
            S0 => ad(4)
        );

    mux_inst_209: MUX2
        port map (
            O => mux_o_209,
            I0 => ram16s_inst_40_dout(3),
            I1 => ram16s_inst_41_dout(3),
            S0 => ad(4)
        );

    mux_inst_210: MUX2
        port map (
            O => mux_o_210,
            I0 => ram16s_inst_42_dout(3),
            I1 => ram16s_inst_43_dout(3),
            S0 => ad(4)
        );

    mux_inst_211: MUX2
        port map (
            O => mux_o_211,
            I0 => ram16s_inst_44_dout(3),
            I1 => ram16s_inst_45_dout(3),
            S0 => ad(4)
        );

    mux_inst_212: MUX2
        port map (
            O => mux_o_212,
            I0 => ram16s_inst_46_dout(3),
            I1 => ram16s_inst_47_dout(3),
            S0 => ad(4)
        );

    mux_inst_213: MUX2
        port map (
            O => mux_o_213,
            I0 => ram16s_inst_48_dout(3),
            I1 => ram16s_inst_49_dout(3),
            S0 => ad(4)
        );

    mux_inst_214: MUX2
        port map (
            O => mux_o_214,
            I0 => ram16s_inst_50_dout(3),
            I1 => ram16s_inst_51_dout(3),
            S0 => ad(4)
        );

    mux_inst_215: MUX2
        port map (
            O => mux_o_215,
            I0 => ram16s_inst_52_dout(3),
            I1 => ram16s_inst_53_dout(3),
            S0 => ad(4)
        );

    mux_inst_216: MUX2
        port map (
            O => mux_o_216,
            I0 => ram16s_inst_54_dout(3),
            I1 => ram16s_inst_55_dout(3),
            S0 => ad(4)
        );

    mux_inst_217: MUX2
        port map (
            O => mux_o_217,
            I0 => ram16s_inst_56_dout(3),
            I1 => ram16s_inst_57_dout(3),
            S0 => ad(4)
        );

    mux_inst_218: MUX2
        port map (
            O => mux_o_218,
            I0 => ram16s_inst_58_dout(3),
            I1 => ram16s_inst_59_dout(3),
            S0 => ad(4)
        );

    mux_inst_219: MUX2
        port map (
            O => mux_o_219,
            I0 => ram16s_inst_60_dout(3),
            I1 => ram16s_inst_61_dout(3),
            S0 => ad(4)
        );

    mux_inst_220: MUX2
        port map (
            O => mux_o_220,
            I0 => ram16s_inst_62_dout(3),
            I1 => ram16s_inst_63_dout(3),
            S0 => ad(4)
        );

    mux_inst_221: MUX2
        port map (
            O => mux_o_221,
            I0 => mux_o_189,
            I1 => mux_o_190,
            S0 => ad(5)
        );

    mux_inst_222: MUX2
        port map (
            O => mux_o_222,
            I0 => mux_o_191,
            I1 => mux_o_192,
            S0 => ad(5)
        );

    mux_inst_223: MUX2
        port map (
            O => mux_o_223,
            I0 => mux_o_193,
            I1 => mux_o_194,
            S0 => ad(5)
        );

    mux_inst_224: MUX2
        port map (
            O => mux_o_224,
            I0 => mux_o_195,
            I1 => mux_o_196,
            S0 => ad(5)
        );

    mux_inst_225: MUX2
        port map (
            O => mux_o_225,
            I0 => mux_o_197,
            I1 => mux_o_198,
            S0 => ad(5)
        );

    mux_inst_226: MUX2
        port map (
            O => mux_o_226,
            I0 => mux_o_199,
            I1 => mux_o_200,
            S0 => ad(5)
        );

    mux_inst_227: MUX2
        port map (
            O => mux_o_227,
            I0 => mux_o_201,
            I1 => mux_o_202,
            S0 => ad(5)
        );

    mux_inst_228: MUX2
        port map (
            O => mux_o_228,
            I0 => mux_o_203,
            I1 => mux_o_204,
            S0 => ad(5)
        );

    mux_inst_229: MUX2
        port map (
            O => mux_o_229,
            I0 => mux_o_205,
            I1 => mux_o_206,
            S0 => ad(5)
        );

    mux_inst_230: MUX2
        port map (
            O => mux_o_230,
            I0 => mux_o_207,
            I1 => mux_o_208,
            S0 => ad(5)
        );

    mux_inst_231: MUX2
        port map (
            O => mux_o_231,
            I0 => mux_o_209,
            I1 => mux_o_210,
            S0 => ad(5)
        );

    mux_inst_232: MUX2
        port map (
            O => mux_o_232,
            I0 => mux_o_211,
            I1 => mux_o_212,
            S0 => ad(5)
        );

    mux_inst_233: MUX2
        port map (
            O => mux_o_233,
            I0 => mux_o_213,
            I1 => mux_o_214,
            S0 => ad(5)
        );

    mux_inst_234: MUX2
        port map (
            O => mux_o_234,
            I0 => mux_o_215,
            I1 => mux_o_216,
            S0 => ad(5)
        );

    mux_inst_235: MUX2
        port map (
            O => mux_o_235,
            I0 => mux_o_217,
            I1 => mux_o_218,
            S0 => ad(5)
        );

    mux_inst_236: MUX2
        port map (
            O => mux_o_236,
            I0 => mux_o_219,
            I1 => mux_o_220,
            S0 => ad(5)
        );

    mux_inst_237: MUX2
        port map (
            O => mux_o_237,
            I0 => mux_o_221,
            I1 => mux_o_222,
            S0 => ad(6)
        );

    mux_inst_238: MUX2
        port map (
            O => mux_o_238,
            I0 => mux_o_223,
            I1 => mux_o_224,
            S0 => ad(6)
        );

    mux_inst_239: MUX2
        port map (
            O => mux_o_239,
            I0 => mux_o_225,
            I1 => mux_o_226,
            S0 => ad(6)
        );

    mux_inst_240: MUX2
        port map (
            O => mux_o_240,
            I0 => mux_o_227,
            I1 => mux_o_228,
            S0 => ad(6)
        );

    mux_inst_241: MUX2
        port map (
            O => mux_o_241,
            I0 => mux_o_229,
            I1 => mux_o_230,
            S0 => ad(6)
        );

    mux_inst_242: MUX2
        port map (
            O => mux_o_242,
            I0 => mux_o_231,
            I1 => mux_o_232,
            S0 => ad(6)
        );

    mux_inst_243: MUX2
        port map (
            O => mux_o_243,
            I0 => mux_o_233,
            I1 => mux_o_234,
            S0 => ad(6)
        );

    mux_inst_244: MUX2
        port map (
            O => mux_o_244,
            I0 => mux_o_235,
            I1 => mux_o_236,
            S0 => ad(6)
        );

    mux_inst_245: MUX2
        port map (
            O => mux_o_245,
            I0 => mux_o_237,
            I1 => mux_o_238,
            S0 => ad(7)
        );

    mux_inst_246: MUX2
        port map (
            O => mux_o_246,
            I0 => mux_o_239,
            I1 => mux_o_240,
            S0 => ad(7)
        );

    mux_inst_247: MUX2
        port map (
            O => mux_o_247,
            I0 => mux_o_241,
            I1 => mux_o_242,
            S0 => ad(7)
        );

    mux_inst_248: MUX2
        port map (
            O => mux_o_248,
            I0 => mux_o_243,
            I1 => mux_o_244,
            S0 => ad(7)
        );

    mux_inst_249: MUX2
        port map (
            O => mux_o_249,
            I0 => mux_o_245,
            I1 => mux_o_246,
            S0 => ad(8)
        );

    mux_inst_250: MUX2
        port map (
            O => mux_o_250,
            I0 => mux_o_247,
            I1 => mux_o_248,
            S0 => ad(8)
        );

    mux_inst_251: MUX2
        port map (
            O => dout(3),
            I0 => mux_o_249,
            I1 => mux_o_250,
            S0 => ad(9)
        );

end Behavioral; --Gowin_RAM16S_color
