--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Mon Nov 06 21:12:23 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_1541_rom is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_1541_rom;

architecture Behavioral of Gowin_pROM_1541_rom is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_RAM_01 => X"808D82101040A0028368F95002D4BD8942706E7A97C8CB40964283284A0A958E",
            INIT_RAM_02 => X"7125BC93888200646411A6592076CB08B11B03894C36F4484036CC2B6C423D03",
            INIT_RAM_03 => X"40E610A19EC0F5A6221331002C7FCF54005B0DB5188460468008D0C067640B77",
            INIT_RAM_04 => X"628C720C0A07E20E40400DD0B33C0064D302133D0A1607FC0828A316888B851F",
            INIT_RAM_05 => X"12217A988830BD34FD68834369265E5A2D15D7F7F4DA23E4BA42942600A62740",
            INIT_RAM_06 => X"2980630BD902C084F23123400499580281801C2D0663038423A2C5A23782B2BA",
            INIT_RAM_07 => X"656868AE51399A2F8B01614DE0688B8368686961B326D8B0C4840A06C19B7065",
            INIT_RAM_08 => X"FE4D0393DD6579678202C80F1816B3F2D8D642DA6D4B48C252D259231E68DD05",
            INIT_RAM_09 => X"AA680B5A8AD15597C480F54D300ECEC64D1E2D9EDB285BFF64961B8C916E4563",
            INIT_RAM_0A => X"9B49C4231101D980430CE5FFA4A3FCCB6ABE8DB6B3B336153DE0B50A7D0D2D5F",
            INIT_RAM_0B => X"E35CDDB224ADF147C23B4851D3832794EF3243EC249998497DD8109F4760489D",
            INIT_RAM_0C => X"E6C4C54804544A0CFAC44CBA0249049898087F3B2B690A2813308CC1842F859C",
            INIT_RAM_0D => X"FDD1E17180EA4D938A44DB04114803030824393149073031E126B20D3525A8F3",
            INIT_RAM_0E => X"211D8209BA602326842B14904A961A28B5DA501E4D2AF87327B8A28FD2D0264E",
            INIT_RAM_0F => X"131849DC8586D5BB5E97E6D3415DC401B47345B2CA686B4871B3018D99242050",
            INIT_RAM_10 => X"189E78887684668C42253CEC808C0002C49AFBD39EA1B0CA2851E680C029A0CB",
            INIT_RAM_11 => X"7B689CB23DB1F0C222DE4332CC99C434F338319439969E1D87031C801C036787",
            INIT_RAM_12 => X"201BC66CB050FB43B81A1B8CC00209EBC475A27AF04898147B9B978809C40099",
            INIT_RAM_13 => X"1E39ED0F871963DE94F96049104F188619F1508B88966C3306A57B67376A96A2",
            INIT_RAM_14 => X"96CFA65ABCFE9BDEB072DE43B7BF43423CFA5BD14AF4C7EA86F0C9DE38858224",
            INIT_RAM_15 => X"2D86F25A90CBDB0140CC4442A91BB44D69701A98BD4D301A4EB784A072F11ED8",
            INIT_RAM_16 => X"E8AF2CB1BCA6096922B25B42C4C0CA0CA044C21E2902EA00BE5128334210658A",
            INIT_RAM_17 => X"28842689BD72C8040473E4E4AF1049259268A045B362C890257A91F0EC65041D",
            INIT_RAM_18 => X"63F39C93A38121C7C4910D9E27E258B504104884080A401848C0303A5859C6AF",
            INIT_RAM_19 => X"751381E8E540DA5462084536825CC17B76412231F8D36E31C11CA1CA2A02BCA2",
            INIT_RAM_1A => X"48D4DD223C308B6D6A9C982D240085865D01367204A72B81D12228022410119E",
            INIT_RAM_1B => X"911A53A3A54E41B2FD272C132CC1668C923720F16A3FA653AD5A6434B4DE75BB",
            INIT_RAM_1C => X"C7938403785F5A2AD30A483074C94058A196BA47913844F69A39C0BA92D31297",
            INIT_RAM_1D => X"4C0859133A9CB808DC15B10B821B006087A0386F213BCE39DE52B0ED8B1432DD",
            INIT_RAM_1E => X"446400CB120536A49E129F4F3831B3D84C68D9A3668D6D27905D311854D2ACE5",
            INIT_RAM_1F => X"E30580C88A392E91A60D5E5A1A6000A839108610AE11159A5E95EF4E39243536",
            INIT_RAM_20 => X"118C6C0230001C5C016245B088D00C717452564699183011698689E3E4066B20",
            INIT_RAM_21 => X"01486CEC1005C00804C8414F90849581FC6F22E737A0E8E73E041F516B8D3320",
            INIT_RAM_22 => X"84772289E4E05E7008211907D9C4EC258312515307887886BEF4E7A86C32832D",
            INIT_RAM_23 => X"98240C58640404834104E998626980BC8375D98CE96B006230557DC36304B4C6",
            INIT_RAM_24 => X"C8460A78038C1CA074C8CC02E42E754D381205231369239508060E1216075B2D",
            INIT_RAM_25 => X"0D45FAAB527628B366C8552A2ADEA6B970E6E2E95AD29AA94D04D62CE16995AA",
            INIT_RAM_26 => X"3C2DA96C36D41440E3700134165386020F6E135FAB446E4010F240A266F510EF",
            INIT_RAM_27 => X"295915A4AD5ED2538A738818CFB28E5620CD301A1A92D0D2D90283DAC91AAC9B",
            INIT_RAM_28 => X"A3493819CEC012BEA54BE76B8CA769C9894EDAA751DB735814161483D4439489",
            INIT_RAM_29 => X"521A992D6E0C4C091C8A45239190714257A5A221C5B8A1C4710A1C4338A21900",
            INIT_RAM_2A => X"04D29E048981A4001045929402030E4180A4120A26B146612B1B1E818A02CA8C",
            INIT_RAM_2B => X"4DA33942956FAFA86DCEDD7395EFAFCDE0CF5ED6919686A824B4E729501FE682",
            INIT_RAM_2C => X"78836F346D9C76F3B7B140CF71030204A0C1A5A232D37AECA4E244DB39B1D529",
            INIT_RAM_2D => X"3E7054D0090CB6D231144DCBDA15346019426B29998119B6CD1B678B2474D676",
            INIT_RAM_2E => X"7B60047888606E8CD1410F92DF978B28E51DC0C646A4FC020F3690239F399145",
            INIT_RAM_2F => X"D01602FBD879136420466FBA7F363E084DFD4FE36324CD4C9A21A0C72B11C6A7",
            INIT_RAM_30 => X"C68A301799A6326EC006D4C6C9B4B2D784134FB353215F0E54C4D27837169888",
            INIT_RAM_31 => X"09709A8D46629DAA5372DF89CA4671B29F61C843CB858D01B1AB4DFA0CD4BE6A",
            INIT_RAM_32 => X"4B04931E0EDD70218A4CD57D7FDDCB4EDA5795494E3052D8F823F06B2468F8A4",
            INIT_RAM_33 => X"624475041454D8962290078A683674B950BEF4CF17281B0549E3C84F8AA2EA8D",
            INIT_RAM_34 => X"766D02B0458924B3EC7D78BAACCF5257B66D0AC3AD438A0E9AAF35BEDBF5C92B",
            INIT_RAM_35 => X"DF55138A68D29230862C01D972F029B325CA41825B73000B0423BAE94F53936E",
            INIT_RAM_36 => X"32F276A3811D1362830898B4CE1221B2C53DE8394E52072C1CA1CA40E538B17F",
            INIT_RAM_37 => X"6D1EA106BB34AD8A01A568FFEBAADDD57382F7F87C01C1FA76E8A7027C877FB8",
            INIT_RAM_38 => X"E2CFD755BBBB99FF911311FFCA2152A33113133113107AB836850E0277C08A24",
            INIT_RAM_39 => X"485739171024C02A166248A5B3AA14A542D24CF1AEB8D7D75DF7BC729E290394",
            INIT_RAM_3A => X"8C9C2D2EE972B18E57541E76BD0D7507B03A7C00D77402EACA0275D7535C7720",
            INIT_RAM_3B => X"997088456F6110C8882081E1FEB6DA80807E96DF3CB9601633B133D80141ACC9",
            INIT_RAM_3C => X"3B013C09F01D0027801F173BF603C50B21B2CAABAABAEA4BC15EDC092C198960",
            INIT_RAM_3D => X"078F67B854820012004DE5CED7E5F020AC00AC53328A8058087F568020A60680",
            INIT_RAM_3E => X"212225757BBBE0DB5AB8614B9ACA540008D4B00001A5694FF7554009EF2E4D29",
            INIT_RAM_3F => X"4FBBBF2092829242A40FA364B3251F037A49BA412D8E932683982C53644666B3"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_01 => X"B800249304BB004808474B4029044A751C0493969504B4080998248000008104",
            INIT_RAM_02 => X"8CD34B690162A111101105B401A2B607A222A40413EDA2C5B509B0C6C1AF60B0",
            INIT_RAM_03 => X"AA455DF2B09520110C162696984108389412D881441105091513736E90D06682",
            INIT_RAM_04 => X"8905A821DF5A8D5AE0CA9B430340A2C18606434050637800114203260521A948",
            INIT_RAM_05 => X"C8DC86A014644861809906285459350290428AA2A290001317B05450C015105B",
            INIT_RAM_06 => X"5A0A960A12649721A7008E1642020250171316A99555294E086800904D080848",
            INIT_RAM_07 => X"DA94C402088471FA88242012509014848985868E6C991304486AB0EC09A6316A",
            INIT_RAM_08 => X"501866A28B5A94003000DA4084084280C80A582108E0044A02408D24DEC91510",
            INIT_RAM_09 => X"5755174244C034142BE28B0407A5250080A12022A289B422924106014F1A010D",
            INIT_RAM_0A => X"045112044B6E80363B090C11651514D04045449504910082CD000021AA828024",
            INIT_RAM_0B => X"56378B4D121B542D1711140088364561426061504116024A0A726D425152B04B",
            INIT_RAM_0C => X"060912EB0A5410884080271104E144004A920A89CA40F2C42089002820107922",
            INIT_RAM_0D => X"A2686140013C646C482230A0090D060050109689088880082081095840202404",
            INIT_RAM_0E => X"552A4D501019B2117302D5266CA210CB29708CD42A4BA601010744217C8D0231",
            INIT_RAM_0F => X"6058A08108D41400141500017A28B6B1A00740301A49284204018CAD122B58A0",
            INIT_RAM_10 => X"B25552E6006AE84653010420A327400010D00C2C555E1AC019AA54481C2C8204",
            INIT_RAM_11 => X"52C4EDA02370208532840090824865161008182084884440512F0A646956D51A",
            INIT_RAM_12 => X"7A9284592D13A6126D04F105961818423CA15E50ADB5A7A3D556C5118D0318C2",
            INIT_RAM_13 => X"20861020A05234508AA10DBC11B40A3031555906CC0459A2C4BD46EA2DD0F528",
            INIT_RAM_14 => X"4E005ED5A0117A94A00284000108CA84A309C4882403CC45001430414004A8DA",
            INIT_RAM_15 => X"D02C5034AD32320350880A0824A462188648463408B248A6D0502404C52EA181",
            INIT_RAM_16 => X"13680127210E00894060228C5B421AA1800095B402C0428C681546D685AEDB34",
            INIT_RAM_17 => X"4A401C206AAC1112FD255B1A126020C211880639A4488460DA80362020803A73",
            INIT_RAM_18 => X"2D421108A895048C524C03609A8DAB43D764590CFEA36A86001102D1A95A9010",
            INIT_RAM_19 => X"A8C5451310B221280965184218B08342222BC006A0115844436214010008A24A",
            INIT_RAM_1A => X"0A1EA0285625A150406B690DA498A00928F7C486D30DC46244C9118C0C604C31",
            INIT_RAM_1B => X"0A28254022A5003120988AF8288001E3D420408F49101CA407AB0D261050A16C",
            INIT_RAM_1C => X"48015B51010804C426D1B5900B1B1887AD4C6A100D15921411520B1404242424",
            INIT_RAM_1D => X"C1AC468805C02404B28370C171D0C20D310C42001A00008000218F1050F5A98B",
            INIT_RAM_1E => X"D609D024C141241004284201080B86BA53850A14081008499002F0E60C006000",
            INIT_RAM_1F => X"00C4623E71004A8D5588B497D55B20034320518C0A630469C0024800024995B1",
            INIT_RAM_20 => X"64E84802202008280008652488B4A820A6D820D2C3085B5A24606008A3BD4A88",
            INIT_RAM_21 => X"20406302082030192059312ADA62D160A8B8C118C0A10208C21341485ECB9901",
            INIT_RAM_22 => X"04212058000640036D688048000029A16281488911451444030B155786B0104A",
            INIT_RAM_23 => X"01C158060269A69829B0046111833589568952111250DE4FA6008AD1204AA030",
            INIT_RAM_24 => X"CC50C023C1BC80002E3C31000000228080014210E30C80894DA08001040A4500",
            INIT_RAM_25 => X"177444863F81540360C4A0CB09DBCDAB6843EB0150D82B00C99A66D95331986C",
            INIT_RAM_26 => X"C0601806E80DEA00202CFB440ED03ABAD55B2015161080C933519E414422E9DE",
            INIT_RAM_27 => X"4200A4040851090022A82483400114043B8ADD83418490D2D105455082710950",
            INIT_RAM_28 => X"18205B408001001460D014044514054880004058000220860800086225B00401",
            INIT_RAM_29 => X"80E0800240409800080002000C99020ED4840DDC008114090205C09101359800",
            INIT_RAM_2A => X"BC23E21A58641F048C2D050802800400181E528010B0360D0161009811F50040",
            INIT_RAM_2B => X"2A140065025054536025888D630114529BB8802000400C07810802164600510F",
            INIT_RAM_2C => X"D31A420BE109A4210D74302230AC2962A015412D80D1514827005F37516C8A28",
            INIT_RAM_2D => X"02100441014000011000D0040063420102090109202CC3A482F84D305203C404",
            INIT_RAM_2E => X"46E814155D03040020008206C188441042E276B93195073041294A6E1022C84D",
            INIT_RAM_2F => X"02240486139034589EDA800A10B4435BD0014213469B60A2A9030C3000036809",
            INIT_RAM_30 => X"34440725221CA1811B5901082A41A108334C046E5A02207B151509CA058480C5",
            INIT_RAM_31 => X"0210412008D92408248520244931804D80544074441258620238121194970945",
            INIT_RAM_32 => X"002030215115101004038A0A8A02901414840280144B8410887A1B4203431362",
            INIT_RAM_33 => X"549A08C220540280913E0115001085500004A4008207F4B89C5D1280141D42ED",
            INIT_RAM_34 => X"800800050024A00556A00C00006362D960001211220004101BD2A81010AA11AA",
            INIT_RAM_35 => X"22210100248008040085503020AA9180021200401005408042C414108AAC4002",
            INIT_RAM_36 => X"E15FED5F7E28004000440212D0D0601C08A20A00042B40012112956908545A28",
            INIT_RAM_37 => X"22945C2014084A15484255410150267FC0016C100BFFBE01EC0416F8227ED577",
            INIT_RAM_38 => X"5168A8A0DDFF11FF911311FFD1122D1008418E08618C10179140E5F8A0BE21FF",
            INIT_RAM_39 => X"400A108203A05ED5628D544021018800354A0428055400A8008150842855A421",
            INIT_RAM_3A => X"1100D0910AA00C000AAA445540EAA21126102A3EA8207155549CAA88AAAA044B",
            INIT_RAM_3B => X"A044307A4A9EAC5402100858CDD2DAD68C22968228100CA14544015236890400",
            INIT_RAM_3C => X"01D48AA41484BA9155C123400010A08A9649B089249209082434407128C8204D",
            INIT_RAM_3D => X"0109248010AA55AAC421408000840D4A0132014957442A0235220C44AB482001",
            INIT_RAM_3E => X"125C4039350DE1AC988D15DC9ADF22244A150149204252A082A058840A040800",
            INIT_RAM_3F => X"E90515448010D22C200012200CA2D440C94019C080408022000000E00041540C"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_RAM_01 => X"043488049009D4001561E32A0646DF9404907460E51ED902D7460361682805AC",
            INIT_RAM_02 => X"33259592821218404049944B2872895128189B231C9248604422C821244B1002",
            INIT_RAM_03 => X"618E58F998C4F001060480262C619C0C73082480400404620048A8A324651BDF",
            INIT_RAM_04 => X"46007328464EC74E30C98D98813030644386A13033100000A269913215988C3C",
            INIT_RAM_05 => X"22272C890E1C381C51E4432364125C6A2E19C7F3E09842EC9921450464444798",
            INIT_RAM_06 => X"398861810962439C612A21034898C00400931E0D8501231E22C7FDD0334792F2",
            INIT_RAM_07 => X"242000502BBD487EC8000304C020410120302120C18390D161208C8341991927",
            INIT_RAM_08 => X"700C50894E14B589741ECF4A950212C6C41C9A5A6C29890820D6C0074378118C",
            INIT_RAM_09 => X"24A44608C285008202F6C534C01CDA0A2408853E583849312590C12413440227",
            INIT_RAM_0A => X"D1024509118997360A41CCB8AC82883B7A7FA01236031211709410086CCCE57E",
            INIT_RAM_0B => X"490A5DB404ADE14787394F04208D63B78C21872014D225177CF9193E754208BC",
            INIT_RAM_0C => X"1ED0C5611670046CEAA004B851703550000075F34FAF0E221710210103520901",
            INIT_RAM_0D => X"F1B0C824A0D5A4B18DC6B983D33462200123525335005A182B05A81D50E08071",
            INIT_RAM_0E => X"21378559E8739B22A32B87B66CD29A40B59999CACF63F44232BAC60EFCDD8E5A",
            INIT_RAM_0F => X"0450619C466CC8F91584E241233CD491A12A64BA5B7D414E1C13042D1C250C62",
            INIT_RAM_10 => X"8814084E92064607130414A8209E4000829E1C41CEE09A0391E8C40844AC9804",
            INIT_RAM_11 => X"522054B030A374E9328C60808D29E106520A19805C884D24091229A418014086",
            INIT_RAM_12 => X"321394683400AA4AA8000BC8104001C2D0E16870B4D80211331144948D100AD2",
            INIT_RAM_13 => X"024A149289091A52049224D000DC48181959584AEA8568AB46946146A2B05300",
            INIT_RAM_14 => X"D45BA46891BE93B424228C60921C952990958BC0361083E248D0701C194B866A",
            INIT_RAM_15 => X"2412700F0CE30B0386A020420D9B7005679148B89DC7D0181E218400F6F09840",
            INIT_RAM_16 => X"88C42491A5242D68129B5A44096212210804C18F00D2E0289E120E24218E8609",
            INIT_RAM_17 => X"31D34F60BC76D84C90D3E5E4A5168A288441060523428114242EB13C6625890B",
            INIT_RAM_18 => X"A3642482425590C64482419226C2409182C54C062C98021102489078C614F23C",
            INIT_RAM_19 => X"FDC0E989612E5A482209861862185A21A88190D1B2580C917A3CA652444610B0",
            INIT_RAM_1A => X"B18866C608AA9824273DAB6C000414824C25A22030C2A23010EB004C2641025A",
            INIT_RAM_1B => X"9221655482DF48A3F36D24BE2890034DD1251275A30BAC66A2E3479011526115",
            INIT_RAM_1C => X"24A785D100C700660348D5C41192253AC590068D9478701A984AE3155464A434",
            INIT_RAM_1D => X"89AC1A10225124048A00A35F36DF574D038613673A19CE38C62134A55358B208",
            INIT_RAM_1E => X"962418EB74602630041AC7052A1D11D20D60C993060C294300CD220A88634729",
            INIT_RAM_1F => X"9150B254D3186CC56699DC1B566BAD705BBD7708A7118BB58B19ECC30BCDC5A6",
            INIT_RAM_20 => X"13CDE8EA36C3041C004143A528FD3C1076D874D4D7521B5B06A229C580F80408",
            INIT_RAM_21 => X"B2164DCC288EE0118570D80EDDA0D1B1FA3D408E5EA00120425225586ECD9B00",
            INIT_RAM_22 => X"52A28410808668401D09D00770100C4DB34D984F0B00B01F871073B82680606A",
            INIT_RAM_23 => X"99C30C4E2768266329B4E4A31260A19851F51B057079DF6376C4FF8800723452",
            INIT_RAM_24 => X"4E0CD2B56119E52436DCD921084AB50641046303624C81864DB4D021860F5F25",
            INIT_RAM_25 => X"BFF29EF5924A73603E3C0BC3640318D1057B33E4A2206430D708A7BBA265C2B0",
            INIT_RAM_26 => X"9845515616A99C280226038403448280ED451913692222CA30D0404544770AA0",
            INIT_RAM_27 => X"230930808CC2D2408EE208106C026D4233CA59931006D8D8DD56059AC21DCD99",
            INIT_RAM_28 => X"8C242D498E44106DA00886220C94254A890A5A25C30B33C614521C63D4A21000",
            INIT_RAM_29 => X"0A08A00C51500E091888442316C1004C8290A66C040014010042C001003A8404",
            INIT_RAM_2A => X"1CB2F20C41619E059045421088082D441687190836591E0606191A1A03100A50",
            INIT_RAM_2B => X"2D833162120C99820F0CCCC718DF734FE0490C4210C2062005B196A89015458E",
            INIT_RAM_2C => X"30DA420A4908642103A318011D631B07428DE8AF300679EA86210E0A3115C613",
            INIT_RAM_2D => X"2A5434DD506C96624223C4CF4B1310021804E12101DB41248292430B0D109424",
            INIT_RAM_2E => X"E143705C5C402E088038EA16891F17412907E60B43A9CE3A4810819318491F46",
            INIT_RAM_2F => X"408C08B2583831066584EC2E56B413309D89CAC34164ECEA8AA3A8C42811C001",
            INIT_RAM_30 => X"C4041115998681000082848250B58100059148135B230C0740D0D26A5796108A",
            INIT_RAM_31 => X"0314098812FBB90877C648E0D022D4B615408560CF97DD6BA4B2049D84871BE7",
            INIT_RAM_32 => X"C8C302FD1E370510BDFAECE46E47BF3DF9CA72BD2C51DE18E932D3E30361B984",
            INIT_RAM_33 => X"160E35C022C4EABAB608220C601940A54288C847DEB80D1D26EB404C688AA6C1",
            INIT_RAM_34 => X"61AD105442A9C096EE577D88C49C6C1A3CA052D68C11C859C2ED10F1247700DB",
            INIT_RAM_35 => X"37700040394E7A544A8012D72F608989159402D4630900954612BE210DD3F098",
            INIT_RAM_36 => X"11DB74E381DCB0D48540AA04CCA0602408378318C21F6319AD7253ED6B4EBBCD",
            INIT_RAM_37 => X"379C60EF8A39C60DCDCE36E9AE7A78784E30F5BC1125C1AC75A0270630874FB8",
            INIT_RAM_38 => X"3AEDCCFCF1F3F1FF911311FFF871954339F29529539F71F01BCC021061800236",
            INIT_RAM_39 => X"824EA50692C0DB6232263C77F3239AD519504679E3BCDD55E4D3A8B5A44FB5AD",
            INIT_RAM_3A => X"640BB4A2814A98BDD1187EF230B4679FF3AD50AB46665A234954511DF110C525",
            INIT_RAM_3B => X"3850383C26A53FA082B08AD8CCF0262A24EB03C65B9769B17701301717100A45",
            INIT_RAM_3C => X"52055822C0A840AB05EC1331B6110501B424000102082140E53AB5780416B847",
            INIT_RAM_3D => X"00466205332A056A0416DCB911982D429542151AD5A8822A0D544B448A862A11",
            INIT_RAM_3E => X"D123B5FE3151E2924E6AD12B0CF15AC001C0305F31CE31B4DCF44082D6E5D4E7",
            INIT_RAM_3F => X"CBEEBD59011600231058510616814C04E9832C04CCD2188AE2D98593098420A2"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE",
            INIT_RAM_01 => X"2F681E0DE2D84052CD4DC00126D65AB44DA63E2027C29B5ED7C6F36B6F6F196B",
            INIT_RAM_02 => X"636CB0B646BA8E67648226D922C4DB9B338C896B15B6D438EEB65D6B6CD9B52B",
            INIT_RAM_03 => X"2DB795A0B3AEE4A223A70B6C644B195D21886D1748E5B86394E589836D2D4B08",
            INIT_RAM_04 => X"E68D2804E645234C2809CD88A136806443402134391500003221B5524C9A8539",
            INIT_RAM_05 => X"2224268C0510941044A643620C36DEC06490908694F38445A16205663C870582",
            INIT_RAM_06 => X"39B2714844A91908FB333B4190831F58D5E8540B063327954262144313A20252",
            INIT_RAM_07 => X"2529289640E58A6B49296404F1288989432129CCF9B37CE628CE090252195E27",
            INIT_RAM_08 => X"9A0D3118182729DAF12AC6000096BB10C440460861382412409214140B726C85",
            INIT_RAM_09 => X"8E88EF008CDEE010E6409218719ED8A4419B8AAA0168D96425B69B69972C2A03",
            INIT_RAM_0A => X"D916871A18DB62B25E2728524420206484802400C88220AC042F011AD1A9822C",
            INIT_RAM_0B => X"E358CA10248DC1275293070DA1A4A93252FCC5DC10716B4409D64C92722A4818",
            INIT_RAM_0C => X"4E886430D4D16C3A41C64C134331199C905875500EA5DE6CA7256B65817CEC9C",
            INIT_RAM_0D => X"6491410D2E40A51E8CE2D31113158E520EA13B33150739312312195406646523",
            INIT_RAM_0E => X"D062A03152222A8000068534DA8430636B17D1150A628019010060E1040D8A08",
            INIT_RAM_0F => X"ED922281A16418C05E46640002610495335E6279337C684040C924099E426098",
            INIT_RAM_10 => X"1E9E238044F8C68F0301000401DDC57CB4D49A9E001CB201A0A172F49522880A",
            INIT_RAM_11 => X"3F69042CA5E0AA9A3084128080806006012138162014B61B050E1708CF5BE233",
            INIT_RAM_12 => X"B27CF61781E6FB13B1DBD94142C8C37B81BDC09EC04D2884799B061CA8B54A9B",
            INIT_RAM_13 => X"1433A90C8400598832C200C4124ED38A34F014C7A83617308C804BC3361A018C",
            INIT_RAM_14 => X"5C045C22045172BCA250841354E9DC5B05A6139118A7821CA600810624A30260",
            INIT_RAM_15 => X"6DA7C35B10FE5ED58ECEC616E09BA44C78A1422C0038A01A94213CBEB0CF5AC0",
            INIT_RAM_16 => X"25E19247109C6D72303B5F96CDD862860A53A21D39104C74387520777218EFDB",
            INIT_RAM_17 => X"51C164C03126554CB0C10CC4C4C81C7182EA226F21C388BA252281582234895D",
            INIT_RAM_18 => X"468D699343602502859764B42D06D9B480F407836589075B969800725A0DA094",
            INIT_RAM_19 => X"E8C20D20C664085A475B2CB0384C230C3260B1A3468325A1E318C42108228498",
            INIT_RAM_1A => X"91C4364624360B0D0CB98320820F1022716C922695E60889064238EB435A16D8",
            INIT_RAM_1B => X"48C80982040941616624309D0989B480D2A62A80C2300438080B432480C831B1",
            INIT_RAM_1C => X"811D6C8128585BCCDC06C1C244500C70C436B2640156E04913942239F10848C2",
            INIT_RAM_1D => X"C58C91A20845F012D815E215841E3E2D80312B631B38C679CE72218C521886DD",
            INIT_RAM_1E => X"145BFA2E00656C96A5CA5260012703B01868D9A346CD043D1012E0E11C086210",
            INIT_RAM_1F => X"48100A0802394011C00C8BC11C03A80F23B81100134BB7061041D9AC33E1D134",
            INIT_RAM_20 => X"3BB09E6002631042BE5A627D002D9041069A2286CE193B1A0610806EC6EA2500",
            INIT_RAM_21 => X"CCC06823832123620C184403DC90C40A0C40122F18A0A0C77244191107C0BA21",
            INIT_RAM_22 => X"80382898504665213C08D00884B542420845910E1D8DD8DD26A780072C802007",
            INIT_RAM_23 => X"BA655926936C062321B1640C2068C409000384489982011C361900C905748D00",
            INIT_RAM_24 => X"CF12C50A9388C202438D8512321102798E98663E264C93126DA2C3CB9C020113",
            INIT_RAM_25 => X"5468B4984A300803203152D310002081411CB3080C0B300BC117730901058400",
            INIT_RAM_26 => X"37A26898933400008478FDD85D02383A676C2A9990526A1605F2FEB27700F48D",
            INIT_RAM_27 => X"58768D6D610842EB0A36DA5BF59B6F7A004C8020639122020EE1D24010227246",
            INIT_RAM_28 => X"BF6D5715ECD7228665D3314CD12649C12D6C94CA9A68480EA8EDA0E82144ED1B",
            INIT_RAM_29 => X"DAD2993F170CDEAD56AF55ABDFEA331681310760CB19B0CC33180CC659B81F16",
            INIT_RAM_2A => X"210C86029A1224608D245BD70AD9EB6CFEFD2FAAA5ED7CEE2940442198E36C8C",
            INIT_RAM_2B => X"80B1ADCBD433662B4A4ED313B5A5CC9A0ACE739C875C80DFB7F7B5B286C06070",
            INIT_RAM_2C => X"30CA4635CD186467176144847D639D0BC28F1F8A2F055256CD42055E19B093F2",
            INIT_RAM_2D => X"0002445600084C0904C9CD85191634074162000B09C91F248D73430824E79474",
            INIT_RAM_2E => X"4BCB61D10BC384FB90100B06830B058E10E6C2DDFD094C28830218BE12D01D42",
            INIT_RAM_2F => X"DA9E10F53794022E6D8EA4EB5E341631D49B6BC74165C9ACA99280B181C76283",
            INIT_RAM_30 => X"72F925661DBC9E2C7CFCD8E6B1B09E9370CE02BE529259EE10CCC9C9254CB4C6",
            INIT_RAM_31 => X"6034424834A06D020D18DA445100CC3680A048470502D4228D2A0DB39464AC89",
            INIT_RAM_32 => X"03EFA1EB55FC26313FED991311B2FF7F6F5EF7FD6E5B5854AA63C6CE204995A0",
            INIT_RAM_33 => X"307A42A694012E8B809480E39937184D1223888953A7E5B40241C409E03400A1",
            INIT_RAM_34 => X"974284DD12E4C4480088802232705C90EAEF0C34489200520288075FFD00C910",
            INIT_RAM_35 => X"62254A4A615EF8DC1B8D769F7F7BA0BE36444694AD7A450DC0A540C6000E23B4",
            INIT_RAM_36 => X"C824BE1DFC2163ACB5C12E3252620C3458A24884210010806316300318C10038",
            INIT_RAM_37 => X"22221C08244A5224025290030190BF99EC893E1126DAFE57BE4E5BF9077BE05F",
            INIT_RAM_38 => X"0408B921FF3333FF911311FF32426FE0B58B58B58A50D94F911BE5E9B2FE65C9",
            INIT_RAM_39 => X"8E1BBD1335C6176D3447B0D6D5892EB45EC00C20080022221181418C60C00C63",
            INIT_RAM_3A => X"E0072538309A343FC4CC2DB18C73128B5FB767B731323899D7D88CC8A0CE1E47",
            INIT_RAM_3B => X"0DE70E05FF39C9A93AB23AF8CD952C1901FF11935FBF17A745E400CDA5209F8D",
            INIT_RAM_3C => X"535C5EEAA7A92B8BDC6B054864F069F86DB6DB33C92492F34349A81242750DF9",
            INIT_RAM_3D => X"5182493C9708DC48DC16FDFF44F984CC37443742B1A64E2E20C112CD8670EA07",
            INIT_RAM_3E => X"F34FB4803381E6000422DE7B4790140F83E0FF9A0A52948183211B82B7EFD5EF",
            INIT_RAM_3F => X"A9502F88B2124127F17B756ED78C2F55B29F34D6A28CBB868BE3F7D766941733"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000001",
            INIT_RAM_01 => X"C81204010890006219604001108153808059544AC82282124141100321604325",
            INIT_RAM_02 => X"600929044106108487628C1A101183A0645152103400014208049B0002120042",
            INIT_RAM_03 => X"300622054008000CC5CF134B484108024A694042B7041653028DC9C048488B5F",
            INIT_RAM_04 => X"D0626D100A6854A14B4C20610001C31A885A40008C20000000A4081016803488",
            INIT_RAM_05 => X"434A46578A2C20AC80888012A8A484B9471D8510018066680A59B685427CE500",
            INIT_RAM_06 => X"8C210A908020025200EC201A2C93996628401D1F0889453C846508A0A545844D",
            INIT_RAM_07 => X"085662693A9590A21B33256DC8662343307C6311F3A741C982119695D2820400",
            INIT_RAM_08 => X"36C0004C0B020005B71451218D042676400102085448C3C933DA0010900CD800",
            INIT_RAM_09 => X"2A128933824A132124A480209114910118903AEB044092200021701214C02084",
            INIT_RAM_0A => X"20602401951005B093436C5000080052501121A124330C630C526110054D6324",
            INIT_RAM_0B => X"C108D88209401AB068C081025048210529092103060916908005862109D98100",
            INIT_RAM_0C => X"1240464EEF282941143B0D40A240A232111022A580310001CB26109002260CB0",
            INIT_RAM_0D => X"60C96E0240694982412AC0B28828416021123320280C2A094880073800961C12",
            INIT_RAM_0E => X"619DAAA0008444CD4CD4080001230E2C94848221B004198CCDD9255452A00608",
            INIT_RAM_0F => X"0038464240820386602861821114446380B300001820C6660C01199C009360CC",
            INIT_RAM_10 => X"4D20C0DD2604612299130C6D319C3601605E1AC29DC194DA5881020128E5144E",
            INIT_RAM_11 => X"32220D05A1B2CC21944221B1409829B2319A0831279CDC9D6603008E82A10C20",
            INIT_RAM_12 => X"05018DA25028496490181B6ECE3858C64C632631909641B03131080B108B3309",
            INIT_RAM_13 => X"313BBC4F12633624CF00C0C822942C5000C3826A390CA2E5C0C8C362E2032035",
            INIT_RAM_14 => X"5697668509659852D43442202000D8A1081AD0A46DB0C0464936000197483466",
            INIT_RAM_15 => X"48C74C9C482A1A57291133443900A90D0859E47204481B4479084341CA1100D9",
            INIT_RAM_16 => X"00620001108624049AB902066DD33A738714991CCC9AC140B9888E5F4916EBD2",
            INIT_RAM_17 => X"6462244000203220040100C8C804D34D583990899020420448445234314E109D",
            INIT_RAM_18 => X"10020241111218346117310100300C216026293409082402212444108190A011",
            INIT_RAM_19 => X"28D84D00E74408509492CB2E53141310CD312008002088089318CB1966450919",
            INIT_RAM_1A => X"2464009184CD1088020999240208123000491A0920020610886E083E85F41680",
            INIT_RAM_1B => X"051A1229111149312144210B445013DC491091F2461DC68D454168A466240310",
            INIT_RAM_1C => X"8C4300DB104F1822C118CD9410DB084918A2130443303420D439E48312131200",
            INIT_RAM_1D => X"8D9CF9F2C2A0A9C98C29B10B0A29196D82921A421A50845094219108D1231448",
            INIT_RAM_1E => X"6C6C18A926619054DA2B58031A11939B64022C0890220425A08B3308C831C18C",
            INIT_RAM_1F => X"5112914DC61825412A2A512A12A233C09223CD935B2DA89AD18C485492490332",
            INIT_RAM_20 => X"33810299849A492300B0240AE602212482C936CC5B320B7B6082081B19308846",
            INIT_RAM_21 => X"633C6499F448B34C439048A2488A5E104901058C113184EC744E9E702AC51B00",
            INIT_RAM_22 => X"38E236102226821364A498A221211A1A9249304B3633630786B0A77065364902",
            INIT_RAM_23 => X"10482806026C32436CB66C870C950A6CA22A2612509534D10080224864415B42",
            INIT_RAM_24 => X"0586D8C0218CB184144C4DA5CE60C0206506624123658584E416993184DA3081",
            INIT_RAM_25 => X"08824100B59115F041C8A4008550214A0C00001C74015FC012C0045658904840",
            INIT_RAM_26 => X"0B208820044004000182050A4089044401C4EEE0103042008048000C88111112",
            INIT_RAM_27 => X"0800402020C000824024160050C8A1080408020808400B0B0088286944004010",
            INIT_RAM_28 => X"4004C0342433390030710CC4330DC36CE4A0544A8A2008166400616412084088",
            INIT_RAM_29 => X"4B034091216048E44A21108940338176C892166608C086058166605900A633F2",
            INIT_RAM_2A => X"D6EC23086DD1119556440943FB6CE536721812E18C840280D0B6406C08182460",
            INIT_RAM_2B => X"810A84E9404000190A140884211100654C6B1CC661D604401242129129BFDF68",
            INIT_RAM_2C => X"4921211E6484921087310840141044381221011A60CC904A7212321B171A08A6",
            INIT_RAM_2D => X"863432C978800030F33248040C2121200312073898091992479924906830DA12",
            INIT_RAM_2E => X"4360582EA220D0066328462240889E71EF07509704B38C9401339D2210244228",
            INIT_RAM_2F => X"855420280407048D6DAD825025C23235F04604AC2269C02D920F040010A12617",
            INIT_RAM_30 => X"02084A0C99844B244504C2C445324B8308029032C040008EB2E2C4104F20CC48",
            INIT_RAM_31 => X"3849C03709C066E50C0091BC27080A0100CA221824C2781E0245C901882C2223",
            INIT_RAM_32 => X"019649AB34849AC92121A802008AA425250840A4A07DC0811584A20018A40042",
            INIT_RAM_33 => X"7CCB86B330D867C9F1044470963408040511B261428007DCC8413F18C60063BD",
            INIT_RAM_34 => X"A41298CF6E79112554AAA911096359742110E118538866703A80431400AA864E",
            INIT_RAM_35 => X"0881B18C6D084F4FE9CDBE14292DCD20D299867384A0984CE6B5545ACBB2DA01",
            INIT_RAM_36 => X"2712714382A8DA1B8CFEE7349488B333E7881A739CEA4E7318C98D48C63552A2",
            INIT_RAM_37 => X"C851C3B514A529D369294D105544776674277142E249C1547141CF04E1071538",
            INIT_RAM_38 => X"D5422088911311FFBBBB99FFD0C8050AB5AB5AB5AB5A5740642A1C268E819C24",
            INIT_RAM_39 => X"270A94E279903440A134D35241110A1034998C8D4556AAAA882452631B352318",
            INIT_RAM_3A => X"DB9600049108932500812589064222494E8500862021301024430888AC890C83",
            INIT_RAM_3B => X"44D84600920040C6DD931E50CC00C321412064CA4A1412234D339F66CFC76C34",
            INIT_RAM_3C => X"C36E4B7259E18DC96E25A252341A311C01B6D8220E38C2034001C20C921844D0",
            INIT_RAM_3D => X"6D80313256436E036E1250A422B2523333D933DB089171E70C08804FF11B799B",
            INIT_RAM_3E => X"81829040371FE16CF38FE008278CCB2065124469A5294A682A886DC252851084",
            INIT_RAM_3F => X"88001616118A010023208439461325B0A92450720220E4B19826120C90301940"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE",
            INIT_RAM_01 => X"8818D6A90BD301C0E1CC6EC066977AB62871555B488F8A6C05549A4C03810B8F",
            INIT_RAM_02 => X"4A09200111A39084853D2E534625CA5126D3D21A9D90016A4AD4D6080A52894F",
            INIT_RAM_03 => X"E427D4A352AC268CD08E7B694DC989446A0F61917766A811BCF12D89494F02A0",
            INIT_RAM_04 => X"F0E8B8D22381D2642730440C24864D36692904860184800011342C993AC25799",
            INIT_RAM_05 => X"2D050B88A186861604A01862EE24C61421069EB6B97228843874A0C56B24842E",
            INIT_RAM_06 => X"04C4216C64927A9819662073A0A10CC18CE5BE49A88991C770B0820E9192C256",
            INIT_RAM_07 => X"0B4C593C94A7D2BB76E2DDC9EF5D337AF04A5AD172A56D60B1015254AEC24490",
            INIT_RAM_08 => X"DDA3C50D2CA308460841AB88425436EBA9442B084F2C42AE567912CC20488AE3",
            INIT_RAM_09 => X"EC08ECAF6B2248D8B4D99D861AD6989C16D26186B0669827000449191625B030",
            INIT_RAM_0A => X"91C1A4C71198704B5C949233B30D3BC48088DA48934CAB2742205AC21D95B12C",
            INIT_RAM_0B => X"6A1A0F15A06061C3CFD3A5A34D0CB3176B903DD91C111A62EC78883371950B18",
            INIT_RAM_0C => X"4572236B4F6B4A4B76490F52CB6F2123147AAA200E739B43882C18C7A848C9A4",
            INIT_RAM_0D => X"64A71D830254361B2C3BF2E86D87B18AA2D81A2586690CAEB4CF7FB146285E5A",
            INIT_RAM_0E => X"C745D54E031113A0A2096EDB81C6629844B7E8826DB2911AA19A1888AB16C108",
            INIT_RAM_0F => X"C385376B314B7015A2989C648E38D9C8C8C49251248235A34692524663926B99",
            INIT_RAM_10 => X"5E820FCD18C1908824C4C6324D564604D5F08D1B2230393464A3243B923F4134",
            INIT_RAM_11 => X"5F4146E1E4CC3382496B4B4D742E9249188CA6A524EB6604A5D8C5BF448BA0D1",
            INIT_RAM_12 => X"12AEDD74774831C796C301EB630D2E6657B36BD9B6044A6559F360D6590C8582",
            INIT_RAM_13 => X"A40A5102E1EE44831D1C36D65C0C380AD57E386F8E047423D7064993668E18E0",
            INIT_RAM_14 => X"79A23142C618C65B99496B4B7CB9604244233891814630C89418D5620831F349",
            INIT_RAM_15 => X"01F160CA46AE4B3924110170B648E4601E6625E6C46E67455121486F9A19027B",
            INIT_RAM_16 => X"38B1249D8431C0681A101FF4E96647665527A8C4147A4B3A88270B2520CBA2C9",
            INIT_RAM_17 => X"80984C9239A63DC4A61DC50504CB0820A0602B6E58B16009210908531132C207",
            INIT_RAM_18 => X"20E31842829BE5E0C416108421C210A4284E2E570024956A21A519121068C894",
            INIT_RAM_19 => X"B968B33D29690859508141050C0B2D891704A46871BE84614DA52C429292C527",
            INIT_RAM_1A => X"01C114070940C229CC0D2E96592848C0396DCB3135348CA5629DAE2C91649612",
            INIT_RAM_1B => X"411610A8DD09D709670C65209765368D20DA0CB535B7699B4F34B5DB4A231935",
            INIT_RAM_1C => X"B94D0564BE1A43461B7292A9452C84220214362114D05B413398D60A9911C0AE",
            INIT_RAM_1D => X"724303074E65FB3C9CCCCF772489439278B4A594ADA52925295A5421A440428D",
            INIT_RAM_1E => X"8B93053D4A972CDF96EF7A518CA268E49508103060C184345D118C2A1710B821",
            INIT_RAM_1F => X"25782F5CD1A7D8C76EF6C2187E6EE88C8EEAA0796CB874A3388459CC36B768CA",
            INIT_RAM_20 => X"AAC73D911DB44513026AF8F68466C5144925492320CCA4849C38BE38C12E5304",
            INIT_RAM_21 => X"05089510DC110E8800AE16F32027282C4C014B2972CD34294BE385CDC73884BF",
            INIT_RAM_22 => X"953960AE2A2B421482552E5112EB4516A5A22DF0B18318342346C88C0E4D14DD",
            INIT_RAM_23 => X"66B6924B2493C99DD248BA29A4C12333A658AD282D228A21691111769DD41358",
            INIT_RAM_24 => X"208922140A5304296312524A208204710A5295BD48B34A5CB279638A51E0C292",
            INIT_RAM_25 => X"00000000000081FF804284048020620482030482814407C5202988000402203F",
            INIT_RAM_26 => X"8455755D02BF3282BA970A12DE68F93B82CD33E0A64B4BB96D60C3260B119000",
            INIT_RAM_27 => X"9C495A7A716842A709349D6F81938631D1FD28D6976936F6F32084DCEC4664F3",
            INIT_RAM_28 => X"32FAFBB8CCE655A22BB325CC9721C959080FF49A9E4C55AB3649BAB45C209A3E",
            INIT_RAM_29 => X"B63CDA26C6CDBD818CC06031992DB687E7E9D56CD19B7EDB368ECDAF9B76BB84",
            INIT_RAM_2A => X"9CB1E4FAC9CF3764850F10856C4906649837648C2F307358DAF4EF8DB5F20CED",
            INIT_RAM_2B => X"1829197086F33775B0463990A535CCC2989C6318C278AD476404232732154589",
            INIT_RAM_2C => X"6DC5B5A11AD6DB5AD1C852B4704A10D304EF23C5112AF26CE742D74C9B3E9947",
            INIT_RAM_2D => X"23195D31AA9E4F10A910E9E51987A69FAA5295E0DB004C5B6846B6DD4146236B",
            INIT_RAM_2E => X"C99ED35CFF54548896863B6FA34B25182182EB596FD30F6523C2153B323338D4",
            INIT_RAM_2F => X"945E41FD7C32EE8C690D8CFEDBEF87B1F19DDB76FA69F9BF741A2F813D79F0C3",
            INIT_RAM_30 => X"6438E495C4379148E236167401879114CE1BF207BED65B03EA2A1C56EFB791F0",
            INIT_RAM_31 => X"96F1E25E8C88A9D41D1293AE47885A01516A2BE1C502914E232BA936FB46E409",
            INIT_RAM_32 => X"37040F2FB5CCB8114049119B9192C046061088C8C7DD25F4B937EACBB2543457",
            INIT_RAM_33 => X"206D99E205B38EA3ACA3CC92183E9B89B732F323812005D0D8693DE99760D69B",
            INIT_RAM_34 => X"BE53F01DC8EB93688F111F336DE6D054F102244887ACC6D21791049E6D11EC60",
            INIT_RAM_35 => X"4CA72B847E111A0DC18F343812399B7226F12CE628733011CD780098D11B9735",
            INIT_RAM_36 => X"142DFA83C1C1973280DC063DB78D2A3DCBEE6A4A529FC94D252A53F9294F3EBA",
            INIT_RAM_37 => X"D90383E0270C6347D8631E3365D4800070E47AD885B7E0867A8D1782867FA83C",
            INIT_RAM_38 => X"3CFB31A9911311FFDDFF11FFC2A445E48F48F48F48F60E0FEC8118161C7F9812",
            INIT_RAM_39 => X"099B195B018BBE48A417828419C7C406F1BD47BA088D1113B9BDCC94A54FE4A5",
            INIT_RAM_3A => X"932C494937137CC666E68235DD6B99209E064526B9BEB4DCCE166EE652ED942F",
            INIT_RAM_3B => X"59D018AB0752128CB8367874CC4D0A655E3C58938C099067C1AAF5C6CCC96889",
            INIT_RAM_3C => X"03CC8E643181D991CCC366DE7F7E68486D249200820820C1EA528AAA96B119CA",
            INIT_RAM_3D => X"C9B060381C564CDE4CE0604E44E32CA00772077622D3A08E5A9994DD852E61B7",
            INIT_RAM_3E => X"3F1601803081E0000000118EB181000FF06A9049646318F9BBA9C99C23026111",
            INIT_RAM_3F => X"F800020458A92CB4CA43387287D74765DE091164B0AFCB66C300A4395725C763"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"C8E3B81D0E11C0C01E40530014874A0C23957044AA04823405855A4601C14B45",
            INIT_RAM_02 => X"420928240E0256A0A1250C1226218269555C1AE2B00041622B84920002128258",
            INIT_RAM_03 => X"8418F5A231AA220AB0CD024D68C3580E439040C1EEE20A520CF15140484BC2AA",
            INIT_RAM_04 => X"B271EE582AE490E05B98A03012016714A8CCF20216037804ABC40A24D3011888",
            INIT_RAM_05 => X"25000442070C028C008808304A34848140828AA280B58440124A0EA07E9AA290",
            INIT_RAM_06 => X"945102D824E92A98CB551233B00000F809B275990AAB410CD0407DF005618045",
            INIT_RAM_07 => X"40040281408690AA9A700A404306A8182501000C48D1840249C5501405022A42",
            INIT_RAM_08 => X"14CAD0182B0210B9702ED7218D852726D4028E001858221180840D23DFF82128",
            INIT_RAM_09 => X"4A84EA33849E333064B48B596104006959919E79E95A90220023F0E284C26EE4",
            INIT_RAM_0A => X"68DF237D81D22B3612654C516D0F14B6D0114DA06DB60C62081D611089696224",
            INIT_RAM_0B => X"4080880309495AB55A51231EF868C9075A02ED528C70E5DC8978C0A26EF9C108",
            INIT_RAM_0C => X"2ED2225F5E430A7B5504C5504A733AAA81C057F7EED60602AF06E71C05400021",
            INIT_RAM_0D => X"205B4B1E103AE802CECB5135DB5CEB3009B5505B5DA853124FB5AF1C4362DD32",
            INIT_RAM_0E => X"C3C4901A011553182A08C5B62082606E4214AA82BB63A41088006C847E8D2E00",
            INIT_RAM_0F => X"9E9376C2E0E62B42082A409204410EA327AA42793A78C6260C49A9B93516418D",
            INIT_RAM_10 => X"0028255460144425DA524849B554EFFCC09008028001149A9881001D09712ED4",
            INIT_RAM_11 => X"10000D20612436B9A6C63135D1124DB420B31221432964B22A42531500000240",
            INIT_RAM_12 => X"3644BF040240BAD7224011408410BB578D2B8695C29621A010382A450C7B10D0",
            INIT_RAM_13 => X"A160105906263C2C4B4AC2093497ED50545530C09A6E04708D98E24070076069",
            INIT_RAM_14 => X"64A004A1021012F6F626C63164689C398116D284F500944069223880A3EBB506",
            INIT_RAM_15 => X"00644B9718B216AA815544306912A1285BDB6EBE400BD85E3D003ED8E88150B1",
            INIT_RAM_16 => X"154092490004C05C302050B46D4F52750161B314B99054182964261E030EC380",
            INIT_RAM_17 => X"752D446828A472A8088D4941408E14510AA6060930E1C2AE0004602E150B005D",
            INIT_RAM_18 => X"765CF271D1E308902105D4210894852808A28F07411345C22E2476100ABCB013",
            INIT_RAM_19 => X"A8826D154A460016969228A0B3443A04235423CB2F30A3C8FA2948200061811B",
            INIT_RAM_1A => X"D54C0B55245F108884081249A4883390086DC40DA01004188A4E12BA01D00550",
            INIT_RAM_1B => X"4442081B30018D61220851166DD8A1508BB0B902C6444695475A6BA622AC0B82",
            INIT_RAM_1C => X"185D289B1280000000300D76209B0851492101684252A6299084040171094874",
            INIT_RAM_1D => X"99997AF5E4A10B39C45926358C1E374D35831342131084508431A1089A292420",
            INIT_RAM_1E => X"26923B320863E459946D6A32131522930842850A142880053400245109084A10",
            INIT_RAM_1F => X"1A2199854E109003806212022007720037724FB96B6BAF16D04158A4976BB1A4",
            INIT_RAM_20 => X"AA9AC55D6F7771CBFE604B17F5BFD9C72CD124CC973313326F1C121C45F03411",
            INIT_RAM_21 => X"A0A0489EC040B49D12128C42950488988952350029351588048AB2308891525F",
            INIT_RAM_22 => X"342538129A84A10378E49AE00D584D4D1A97B0DE288B88AC0200A0004526B36B",
            INIT_RAM_23 => X"32E32D249269B4FB4D32690B16B1AE6CA2688AD0D911BE66348022D369E1328C",
            INIT_RAM_24 => X"CB24C1017109C206058989B0100100410B88620A3669350EE934C2C18E4F3893",
            INIT_RAM_25 => X"BEEFF7BDF7DF3F007FFCBFFBFFD043FB7DFFFBBCFE45F818DFC037FFF8FDCBC0",
            INIT_RAM_26 => X"AC421084250804004C04F6D2C7833C7EA0E066A8083444DF344A2C0CA90017F7",
            INIT_RAM_27 => X"10244C4C40C000B8462456C7E0C14421D5D80AE620193ADADF622658D5045230",
            INIT_RAM_28 => X"1E48DE308403AF001E310EC43F0FC2CC8004942A8E0454D468496D4526A08C13",
            INIT_RAM_29 => X"D391CCC35266DBC8884020110F739B6EC923010260CDA66D9B2466CA0DBC1F40",
            INIT_RAM_2A => X"FFB0E3ECFFE117D457054003FEED04369C043F840DF82CEEF06264DCD9F94466",
            INIT_RAM_2B => X"E90A10C00351151B6014A884000100580A0825086E6805D04000020BBF376F8C",
            INIT_RAM_2C => X"591B630A4D8CB63185220C6038435801542B13014988D05866005E12038A88F6",
            INIT_RAM_2D => X"842634DE41CC4E0884CDC8C406022A6F62141677815A0136C293659448009E36",
            INIT_RAM_2E => X"424DF3D7A8D35479835CEA268109068610034611053BC53CC18005A291C29F4A",
            INIT_RAM_2F => X"845481D01B9274294DA9A4AA5E76A2B5B4994B4B6A4958B5929B8C8091654455",
            INIT_RAM_30 => X"001B424E4405C50003A40A145502C5000B829082D6D24902B26A44534D6DF09A",
            INIT_RAM_31 => X"5355C07A78E8A344140891FC5728C0A58142A2CB64D27C4E9E768911294C6281",
            INIT_RAM_32 => X"0165014328E09CE00004888A880880840001088085EBEEB5ED7742469AE19562",
            INIT_RAM_33 => X"0A016016109B0350F11580825107084022022BBC081016BE0B1DA934A0554A48",
            INIT_RAM_34 => X"771CDC067039D64916222C00127A140888460DA78C0F3829520B34570000C3D5",
            INIT_RAM_35 => X"2203D1420C010F8670C1D810802EC93880D5604200B9FB4866A0AA040000F381",
            INIT_RAM_36 => X"E91FE1433E28B397E9674B0486EBBC006000A494A52312964A4CA46252905800",
            INIT_RAM_37 => X"22705C3D11E318706318C140100000006849610323FF9F546146567D21061533",
            INIT_RAM_38 => X"41608800911311FFF1F3F1FFE08E670ED4AD4AD4AD48C140113805E1820065E4",
            INIT_RAM_39 => X"B30210420F540544A155AA200D0060002A99810D44468888000817294991894A",
            INIT_RAM_3A => X"A29500041080414422ABC61D47DA8A718514211DA803EC55778CAAAAF6A0D64E",
            INIT_RAM_3B => X"097F0842001080E7EC136C50CDB2AF3C1A35358A884094630122197DAF039E20",
            INIT_RAM_3C => X"80760BB05EC00EC176058218363038630536D910410450300006E08E0C1C0961",
            INIT_RAM_3D => X"C054321ED54E7607E600420722A8DA7F21DF219B99E23D430C200046D223B01D",
            INIT_RAM_3E => X"65C70180302143FFFFFC7FFE251EFE1AC0320AFF8718C6000000FCC042102010",
            INIT_RAM_3F => X"E8002EED2604D2607801603001120580D2A09C601024C13281C4001813809A51"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_01 => X"E7CBA2B0EC4B3D52BB6DB37F52D0F79CA7353D3ECA1E5B4883D2A12842084286",
            INIT_RAM_02 => X"29649D93DC974EA6A5BBE8C976FD19EB554F49C938B6812AE7324B6B5AC9B171",
            INIT_RAM_03 => X"C18B66032A04D54AA7EF79252520C45F299B2DEBEEE59A52B67CF0EB2525D9FF",
            INIT_RAM_04 => X"76E29F1CE76CD6EC3B89ADB9B33563744BCC93343737078289C5AB26CB1B98B4",
            INIT_RAM_05 => X"696F7C5BAF3CB4B8F7E6D37664125E752FBF2F2D0088EFEDD93FAEA53FFAE63A",
            INIT_RAM_06 => X"B59161DB5B66D1CA59552959BCBBDD7FAC9B1B1EAAABC7A2A7C7E9B233E737F5",
            INIT_RAM_07 => X"6D6D6BE5F7FFCA57DA3B534D2B6FAB5B777B7B5DFBF7E1A1EAD54F53A9997266",
            INIT_RAM_08 => X"FCC7455967273973A774933F399637E4997EDCDED933FBB935C6DD30004AEB8D",
            INIT_RAM_09 => X"666E6733DCDB6336E2764F6DB30E4EE5598B9F7DF5304B136D9673CA928E6CE2",
            INIT_RAM_0A => X"A95CAF33B4C93DA44F61E9E9E9CF9C9B7EFFEDA6B7B36C73FDBB638A4CECCFFA",
            INIT_RAM_0B => X"F90E57BF24243870D02BAE39D96746B0B58F43BA9669CCD374A2CA9D0AB14A94",
            INIT_RAM_0C => X"74C0CD2D7AAB4734AA154EABE9399AAA958AFD7001AD8C36AD2FCE58AE6EC5BC",
            INIT_RAM_0D => X"D1F9EF795EFF69BBC367EB269A6D4772AFB639326D0F3331C9B31F3FF5B39CF3",
            INIT_RAM_0E => X"F5FBCA99FAF7757DEEF3C1B648377EEFBDAADBBCF7647DD6EFFFE61FFCF924DE",
            INIT_RAM_0F => X"591827DAEDDEF3B62DABE5926BBEF6B3A6776DA6D34CE63E7CB78D9D135F7ADD",
            INIT_RAM_10 => X"0AA8BADD66CCE3BCDA1F39CDB19B7EFD159A97DBCAB4AC9B7BFB97689C7F34CF",
            INIT_RAM_11 => X"7C32F91110F3C673A6DEF331CCF1CDB4E6B331BD3B1EDE9DA63B11E472298B9C",
            INIT_RAM_12 => X"80E3DF713D067157159B4AC9869959E7FCF3FE79FC462F373E39CB9D85E6185B",
            INIT_RAM_13 => X"3D39FD4F163B77AC4D78CC7D32459D42A9EFAACC5F6E7173D2B8A1EC73EBE6A9",
            INIT_RAM_14 => X"FE5FF69B35EFD9DEF676DEF2A2959B7334BBD9374DF6C3FEEDE3F99ABBE9323C",
            INIT_RAM_15 => X"6D032E8C5C7D094209555446BD09CDC52E31FCFFB76E314CBD2943C5EA5B804A",
            INIT_RAM_16 => X"98CD6DB49CF6082EB2920C46EDB31B7591465B88EDD2984891C0AC7F6B9CEF9B",
            INIT_RAM_17 => X"44AE78C99DD3AAA49C76E4ECEF74CF3CAA77AC67B366D2966D7E6364DD6B9A86",
            INIT_RAM_18 => X"5279CB5397B32EF6EC93159564D254B5AE62A7132CBB4399BCB5746ADCB866FF",
            INIT_RAM_19 => X"578BEC98E73CDECE52C9E79DD15ED26BCF5597293CB2AF2BD21CE7FEE6E7B4F9",
            INIT_RAM_1A => X"64DCDD93BC5D0AED6E34F36DA68773925F24E62D94A3DEF9CFEF707E57F2938E",
            INIT_RAM_1B => X"B7B5FF6B13DFD9B7D3672CF36CD927DF8BB2B9BE673BBC56AAFA69B462ACC39F",
            INIT_RAM_1C => X"ED5607DB385F5B76DBDE792677D3673F0D921D477F607666C77FD3C726FEBEA3",
            INIT_RAM_1D => X"8D0C79F3A651C5B5CAB8F2DD6DBBDB6937AF3A6F733BDE39CE73BCE79BE1B240",
            INIT_RAM_1E => X"846D58FFF6E5DABEAB9EF54E7333A17B1F3A74E9D3A76737B1DFB3FFD8FFC9FF",
            INIT_RAM_1F => X"FBE3F9FDF7796CEDE781C899D67B33ECBB33EF8A861B1DFBDFFC84DEFB6DB127",
            INIT_RAM_20 => X"336F739DFDBE555F7E8ACDCEF7F6ED557491F68E9A3B321B69E6F1B31D3AB113",
            INIT_RAM_21 => X"7FBECFDDF35DF13F5BF07CEF90EE8BFBFD7FF3E5E731E4EF3C8E9E3B66CC9B21",
            INIT_RAM_22 => X"BCFF3EB1F3ECDFF768E798EFFCC8191DFBDA3B93763A63B6A5F6F2AD2B26D347",
            INIT_RAM_23 => X"99E638DC6E49B4DB4D23E9E33A74ED5955F4BBCAF87BBECFE4DDFF9B606562F6",
            INIT_RAM_24 => X"A9BE9FFFF33DBFEE72FCFD33BEFFFF5C6196E737F36933B869369A7B94FE7EED",
            INIT_RAM_25 => X"A2A814A51450028000A14A01400A95000004814140AA08228016400A01401440",
            INIT_RAM_26 => X"99EFBBEC97DDBEFAC70E0F42DE8B3C7ED8E7552E77746EC930EA5E2AA8DDBA14",
            INIT_RAM_27 => X"735B79C9CD8EF6595CF28C9BC5C38A5237837BBA7B56D393910EAFF1877FEDDF",
            INIT_RAM_28 => X"B26CBA298AC18F79D4AAAAAAAAAAAACC090ECFD5514B238C78B6F8C7E7EE39B2",
            INIT_RAM_29 => X"9BB9CC86676698C91888442319199A7ECBB3923A6DCD36699A27E68B0D27B140",
            INIT_RAM_2A => X"EF4557F67E26ABF5DF6F9296FEFC4C7E383A74882B316668F6B61EFCD2F80EE6",
            INIT_RAM_2B => X"44A93162972AAEB3454E7FD29CBFEEDFDA5F7FDEEFFEAA20049CA6363FA8CA35",
            INIT_RAM_2C => X"38BB673F699C767392F17CE7712849C39CA4E105508AABA8AB02CB0F63955545",
            INIT_RAM_2D => X"FCE6669B5BCDB6FEEBBECDDFD73736631BD3E6379B09DDB6CFDA638B67F6DE66",
            INIT_RAM_2E => X"A1EE9BAF01B0AAF75769C766DBBEBFEFBDA7AC4FEFA3CB24DB12949989939A68",
            INIT_RAM_2F => X"D05700CCE06E32AD6DADFA9739761535BF44E72B6165A57FB36FFC4D7830C292",
            INIT_RAM_30 => X"E76F272F9DB2CF6EE616D2E765BDCFD7C63BC825C925160D62DAFAB22E92ED8C",
            INIT_RAM_31 => X"3239DBB665FF3AC5F7D6D3BDE76E73933E6BAAAAFFFFFFDFF9558D2B180AB32B",
            INIT_RAM_32 => X"ABAE03962B8A92E1484B55575555C9CA4A5298898A7FE4495F572FA93EE4E8CE",
            INIT_RAM_33 => X"2A65555685DB4E53A2AA2A28A02C5CA150A872AA92282FFD58AB2974CAA2E64C",
            INIT_RAM_34 => X"7455DC9DF4E91492AE555CAAA4C738CA5554A94A052AAAA89B5550AC49558EC5",
            INIT_RAM_35 => X"5555CB885C531B9CF38FF4B9827F99A285D94CC209E3DB49CC6200AD55599225",
            INIT_RAM_36 => X"1A0058A2C1559233E8CF463CCECA7D3AF5D57DAD6B5735AED6AD6AE6B5AAB975",
            INIT_RAM_37 => X"5568A172ABD6B56AE6B5AAAAABAA8000729A58AB400160A058B2858340858A2C",
            INIT_RAM_38 => X"AAE57555911311FFFF3333FF8EA94429CF5CF5CF5CF5A2802AB40A034500CA00",
            INIT_RAM_39 => X"275731442B968C6AB557C20493A29485F5D94A5CAAAE55555552AF5AD5AB9AD6",
            INIT_RAM_3A => X"CAAE252AB942A88C55D7483BBEC775529624532E756572BAEC945D5555D54423",
            INIT_RAM_3B => X"405F42A5232949CFF83378F0CC008373546C74D71CC17C9622722BBCEF6BBCA1",
            INIT_RAM_3C => X"13FC9FE4BF895F93FC4B173976D179DD25A49332CB2CB272A948CA9E54F90059",
            INIT_RAM_3D => X"55A27931BE4AFC4BFCA4E60C55F2AE7F277F27733988BD4E585552CDB287E2BF",
            INIT_RAM_3E => X"B3DC24003001800000005FFE71A001056062156996B5AD5557557F94A7304531",
            INIT_RAM_3F => X"B8003BF5B1A6D362C00BB1709393CF81BA2131E0ACA6C3B003B424B852053A53"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_1541_rom
