--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.9 Beta-4 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Sun Dec 31 18:51:07 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_1541_8k_rom is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(12 downto 0)
    );
end Gowin_pROM_1541_8k_rom;

architecture Behavioral of Gowin_pROM_1541_8k_rom is

    signal prom_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= prom_inst_0_DO_o(1 downto 0) ;
    prom_inst_0_dout_w(29 downto 0) <= prom_inst_0_DO_o(31 downto 2) ;
    prom_inst_1_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= prom_inst_1_DO_o(1 downto 0) ;
    prom_inst_1_dout_w(29 downto 0) <= prom_inst_1_DO_o(31 downto 2) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    prom_inst_3_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= prom_inst_3_DO_o(1 downto 0) ;
    prom_inst_3_dout_w(29 downto 0) <= prom_inst_3_DO_o(31 downto 2) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"8042CC0153301F011100560617304D8071018270149041500C04218C1CF0083C",
            INIT_RAM_01 => X"30E0558011489D844522A4535169D46115858D047472008E248C09900088D93B",
            INIT_RAM_02 => X"048C96E1920594E21094C20C3899F0D10540014C107CD11CC4134CA451178192",
            INIT_RAM_03 => X"4B0148C41621DBD441601D3DC416361BD445201BC888056D0474137482329A04",
            INIT_RAM_04 => X"7864594E4253070D103899F0D14350C0900441C925A020814807114885911480",
            INIT_RAM_05 => X"01C7058859181601281058C7058636F5141418D3DC405D886F51C1601BC08F32",
            INIT_RAM_06 => X"44146852082A045208A05347025853080517074211634604D411C12C80116816",
            INIT_RAM_07 => X"378D55A5108A491C0088343042151C9148A01452161C11484D9A148998681489",
            INIT_RAM_08 => X"544640012344D3B90D00160001051047676DD5855019DD993216451E22344E01",
            INIT_RAM_09 => X"058045051D5888F330424756A0E07416110763367008409148220302455D166A",
            INIT_RAM_0A => X"26675099998C0A1C819C0038141434401324491610A99A91A99A916044B3C181",
            INIT_RAM_0B => X"2119182748B3C9031494430F30415070F1C85058603945C99D004CC266549991",
            INIT_RAM_0C => X"6011414756223CCC12507C7011414D0452505801324191E10211912111121191",
            INIT_RAM_0D => X"C998C0A3C8CD9C00381F30004CC192245842826682468266824644112CF07041",
            INIT_RAM_0E => X"A68114E141C45131146A46159A1D99104345C9D004CC26425499C91266277099",
            INIT_RAM_0F => X"549110007604C00440937254910254766AC106428D593766460190229A041188",
            INIT_RAM_10 => X"0050920050741305019044114400415420190608C00701505200133003B14D10",
            INIT_RAM_11 => X"852188A303210841655024091A1C31948118053374423081000504411694C012",
            INIT_RAM_12 => X"08886088950050951215A55A2053000855C530C016A3CA0CB14A383215A56194",
            INIT_RAM_13 => X"15A5487345C1412254040510614314219620A54232150885C01533506537514A",
            INIT_RAM_14 => X"450AC95DD28E0D1209041818A18462624250C9E314088BD61CD96161500191A2",
            INIT_RAM_15 => X"6299C1434198590541934612A509850434041424A85509050059154DC904594B",
            INIT_RAM_16 => X"90D5A55837410C4179A62D1B2564456616D4DA404094541A414344444042514C",
            INIT_RAM_17 => X"241D5420D3444C015C0514561556A9349C4428407027459100101D7091890708",
            INIT_RAM_18 => X"449143653402D1E405882C1C0065265C81CD9C003845051C14022D80684D9433",
            INIT_RAM_19 => X"99140071C104D10399140147041A9187668664502704182645005C0021819996",
            INIT_RAM_1A => X"89062C485186227661214B4449128366369DB446D5594650C60C104500CC1040",
            INIT_RAM_1B => X"D2045F36A748916C04495155746695C100101DA0917224182143440712361A44",
            INIT_RAM_1C => X"445000704199916001C10664458007041264540070411DCF0455451251C1BCA9",
            INIT_RAM_1D => X"6499199D15CA55011699114001C10464A9D204548A7489153099915001C10664",
            INIT_RAM_1E => X"0D10659440155964155944155964155944455659C599A598416C3468C3A1A852",
            INIT_RAM_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF64",
            INIT_RAM_20 => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_21 => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050",
            INIT_RAM_25 => X"FEFEFAFA54545050FEFEFAFAFEFEFAFAFEFEFAFA54545050FEFEFAFAFEFEFAFA",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555555555555555555555555555555",
            INIT_RAM_29 => X"AAAAAAAAFFFFFFFFAAAAAAAAAAAAAAAA55555555555555550000000000000000",
            INIT_RAM_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2C => X"AAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAA5555555555555555",
            INIT_RAM_2D => X"AAAAAAAAFFFFFFFFFFFFFFFF55555555FFFFFFFFFFFFFFFFFFFFFFFF55555555",
            INIT_RAM_2E => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_2F => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_30 => X"000000000000FFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFDE7D7F2DA884",
            INIT_RAM_31 => X"FFFF00000000FFFF000000000000FFFF000000000000FFFF00000000FFFFFFFF",
            INIT_RAM_32 => X"C303030F0203FFFFC303030F0103FFFFC303030F0203FFFFC303030F0203FFFF",
            INIT_RAM_33 => X"C303030F0003FFFFC303030F0003FFFFC303030F0203FFFFC303030F0003FFFF",
            INIT_RAM_34 => X"555500000000FFFF555500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_35 => X"FFFFAAAA5555FFFFFFFFAAAA5555FFFFFFFFAAAAFFFFFFFFFFFFAAAAFFFFFFFF",
            INIT_RAM_36 => X"000F000F000F000F000F000F000F000F0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF",
            INIT_RAM_37 => X"F00FF00FF00FF00F000F000F000F000F000F000F000F000FFFFFFFFFFFFFFFFF",
            INIT_RAM_38 => X"E7E7EFEF4343FFFFE7E7EFEF4343FFFFE7E7EFEF4343FFFFE7E7EFEF4343FFFF",
            INIT_RAM_39 => X"E7E7EFEF4343FFFFE7E7EFEF4343FFFFE7E7EFEF4343FFFFE7E7EFEF4343FFFF",
            INIT_RAM_3A => X"FF5FFF5FFF5FFF5FAA0FAA0FAA0FAA0F5F0F5F0F5F0F5F0FFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFF87E943A50B61C72D83E94ECECECE8A888884464646020202CECECE8A8A8A8",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3F => X"03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"5F6D7082530073C720E0972832008B81D00170607420F3ED33D38EF7C70C78CB",
            INIT_RAM_01 => X"C073CA52CCEC498E33B2A33A63549CE525B3C98D5B3B0144164307A41088B21C",
            INIT_RAM_02 => X"8AC554554B25405B132430F01C7A20722D9041302CCF1048D422C094F51D0710",
            INIT_RAM_03 => X"D42CEC4ECF139894ECF139890ECF243490F3B034C8ACB34EFCBBFCFACB325960",
            INIT_RAM_04 => X"555254054C90C1CB281C7A20724D8302CB3CB2020E70B2CCEC4C3CEC0D43CEC0",
            INIT_RAM_05 => X"130D33C0D434CF035C933C4F334F262530CD3C9890D339C0D2434CF034C94415",
            INIT_RAM_06 => X"8F14AB3B0C1D173B143CB2CB0FEBBC244B2225B2D2E2CA08B029428F1CF298CF",
            INIT_RAM_07 => X"2C45CA572ACA09943EC805273B26309CECA8273B263C9CEC856ACEC998EACEC9",
            INIT_RAM_08 => X"4485904122C8B1C53202CD33C9E722655562558964915151023D4754322C8782",
            INIT_RAM_09 => X"3E501CC73D195D3C144CB9C87073F8F9C5B056145800486CEC5140C1CB7FDFE8",
            INIT_RAM_0A => X"A6707299C15415575914141014CA164407642C0192DC8DC8DC4DC06E40310182",
            INIT_RAM_0B => X"155C04F154310D4373DCE143C0B3AE123C4423E58255B20991101DCA671699C5",
            INIT_RAM_0C => X"940731CF46574F051371CF10F24C8B3CB371E4407725C0D92155801558015540",
            INIT_RAM_0D => X"4C154155758514141016DB101D80983006CB432363234313630130900C40408F",
            INIT_RAM_0E => X"96580A41738A52C558EA16356A8141054DB2091101D4A66316990C5A66304299",
            INIT_RAM_0F => X"C8B28E3BE92F88CAF020D264B20266556AC23EC2019094546707000259602900",
            INIT_RAM_10 => X"2320A32328DA3AC5A328E392848DA3ECA2328D2008D923E8E12369E238C2632B",
            INIT_RAM_11 => X"48C648BF8B226489985929816BC0926248E4C123B96900B212328EA38CE888E0",
            INIT_RAM_12 => X"A41A90BC19D09C22B0693A26929C8B21A4C9C0EC96930BC89E8BC8A0693A0662",
            INIT_RAM_13 => X"693A249D68CA7410971989C09E74088262923A77307BE018CC61004286386041",
            INIT_RAM_14 => X"C801421E51834DD0821C20F4020CA09091B70AAC0B368BF42CA0C0879D4A7250",
            INIT_RAM_15 => X"30BA8E00C328EAF48720D8303A021C1A090809185042421C124A93BA020E4BE0",
            INIT_RAM_16 => X"B015A4AC8FA8C0891E78032518588599283C20D282AC6020C0A14A48B18281A3",
            INIT_RAM_17 => X"047D11E018CA388CA449BC89A24AA5CB60552454F20E8368E3BEFABCB2420B20",
            INIT_RAM_18 => X"169500C00410B2D4C9430CC441C3253046C51414101CC73C24C70E83AAC10030",
            INIT_RAM_19 => X"998E3CE28BCA125C998E358E2F2A858C5AA26638D22F28A6638C309728E39994",
            INIT_RAM_1A => X"C54DB0EC520EB0445BB1B2C4883033B4161E2D4A1922C8B8CC88BCA38F78BCA5",
            INIT_RAM_1B => X"EA423CCAA7A988F71C8360D854569788E3BEFABCB2E108208248CA253B15314E",
            INIT_RAM_1C => X"22388DA2F29948F2368BCA642388DA2F2A623C8DA2F205C4061C872A1BC973A9",
            INIT_RAM_1D => X"5654199581CA500F219908E2368BCA10A9EA6230AA7A948C329988C2368BCA66",
            INIT_RAM_1E => X"CB21C662CA166621166620166613166602859988C9296584A8F72CBF0A414402",
            INIT_RAM_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA1",
            INIT_RAM_20 => X"FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050",
            INIT_RAM_21 => X"FEFEFAFA54545050FEFEFAFAFEFEFAFAFEFEFAFA54545050FEFEFAFAFEFEFAFA",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555555555555555555555555555555",
            INIT_RAM_25 => X"AAAAAAAAFFFFFFFFAAAAAAAAAAAAAAAA55555555555555550000000000000000",
            INIT_RAM_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_28 => X"AAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAA5555555555555555",
            INIT_RAM_29 => X"AAAAAAAAFFFFFFFFFFFFFFFF55555555FFFFFFFFFFFFFFFFFFFFFFFF55555555",
            INIT_RAM_2A => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_2B => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_2F => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_30 => X"000000000000FFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFDAFB94EE6B44",
            INIT_RAM_31 => X"FFFF00000000FFFF000000000000FFFF000000000000FFFF00000000FFFFFFFF",
            INIT_RAM_32 => X"C303030F0003FFFFC303030F0203FFFFC303030F0303FFFFC303030F0303FFFF",
            INIT_RAM_33 => X"C303030F0003FFFFC303030F0003FFFFC303030F0003FFFFC303030F0303FFFF",
            INIT_RAM_34 => X"55555555FFFFFFFF00000000AAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_35 => X"FFFFFFFFFFFFFFFFAAAAAAAAAAAAFFFF55555555FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_36 => X"000F000F000F000F000F000F000F000F0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFF",
            INIT_RAM_37 => X"F00FF00FF00FF00F000F000F000F000F000F000F000F000FFFFFFFFFFFFFFFFF",
            INIT_RAM_38 => X"FFAB5F0F5F0BFFFFFFAB5F0F5F0BFFFFFFAB5F0F5F0BFFFFFFAB5F0F5F0BFFFF",
            INIT_RAM_39 => X"FFAB5F0F5F0BFFFFFFAB5F0F5F0BFFFFFFAB5F0F5F0BFFFFFFAB5F0F5F0BFFFF",
            INIT_RAM_3A => X"E44FE44FE44FE44FE44FE44FE44FE44FEFEFEFEFEFEFEFEFFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFF9B6546103DCFA8B657210FFEEDDCCFFEDCFEDFECFDCECDFCAB9A89B8AB9A8",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3F => X"03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"A48243142B8C8D08228608502A87021226F8AE9C814090928928A28824928920",
            INIT_RAM_01 => X"0C0049B414BD14CC52F6852D33654CE4A412D4CD092F4A2B9AB9806AA6D01200",
            INIT_RAM_02 => X"C9D662447F44726F60219A010006B80200AA9B0164B0D8AAC1C0AD04B52C88A9",
            INIT_RAM_03 => X"DB443DCF4371634CF4371634CF4353334CD0F737ED3DD02E4019243BDF641041",
            INIT_RAM_04 => X"911C472680866800210006B80280A0302007AA1409B2F7D43DC7343DC5B343DC",
            INIT_RAM_05 => X"71CD52DC5B394B7369352DCF52C758D3314B1D634CD524DCCD3394B737EE2899",
            INIT_RAM_06 => X"CE62A12F6900E12F62C0000B643CD042802A818C6020097029C2B66C901A614B",
            INIT_RAM_07 => X"0CA4DD137BD014410FD9C1612F533984BDA7612F533D84BD18284BD44CEA4BD4",
            INIT_RAM_08 => X"B0B0AA9B4040300A028B4BD2149069111A02A80ABE4A4646B424C972A4078236",
            INIT_RAM_09 => X"0DA6CDF378ECC8D0E680A54AB400783616059841BA2D0014BD890E60083F0FE2",
            INIT_RAM_0A => X"33259CCC96E8B32CEC68B0AEE80943B0B2B3C8FE24A83A83A83A8F933CBA2E3A",
            INIT_RAM_0B => X"ECC9E824B0BA2A9A378DF66D0592E288D22300588F88A21CC6C2CA133258CC96",
            INIT_RAM_0C => X"69B37CDE3B3234398F02B4881A8080078F029B0B2A4C9EA14ECC1EECC1EECC1E",
            INIT_RAM_0D => X"596E8B320E9068B0AEEB2CC2CA1DE163F852A60EA60EB60EB63E81CF2E8B9E83",
            INIT_RAM_0E => X"0410492931CE4A344CE8D334283434FE80A21C6C2CA1331658CC99633065ACCC",
            INIT_RAM_0F => X"080249240BD294992F40BF3802891111A0120EFA104F11919248F2B4104124AD",
            INIT_RAM_10 => X"D22536D224392920500492C2F74890ED09004B49F48890E4B4D2293D24079024",
            INIT_RAM_11 => X"680AABA0A661E63E742DE1A02A1A75D2682AF69C0899B42BCD22401240FD74BE",
            INIT_RAM_12 => X"6A28942DF91290D26417359CAA91A4705DA91232CA0D6A2A822A1E64173589D2",
            INIT_RAM_13 => X"1735AAB309AE46841851A92A92449675D8AA3644AC6B310DA7069CACBCC08DA2",
            INIT_RAM_14 => X"388A2E02E00A1C62340810A26200A504852414A05252D3D221808C0E916565CC",
            INIT_RAM_15 => X"2882109000618910806228682A703A5048514841469A140A4A9E26AA340C9AC0",
            INIT_RAM_16 => X"AE0030AA43B02D427DFC80E8A801801A602900B62F2FC1C097072303871F3D08",
            INIT_RAM_17 => X"E0A8E11204092D48AED56267994A082AA3258925892288E49249028002D40CC2",
            INIT_RAM_18 => X"58C4B237D8B452E8080A2E22F23C70E652B068B0AECDF375A8082210E230F2B8",
            INIT_RAM_19 => X"CC412C73F49A4AC3CC4124CFD26A34CD0A0F31048FD26773104BE6384412CC9B",
            INIT_RAM_1A => X"D8C4ACFD80CEF6110AF54146A0602BAC6E022C220C2300EF626F49904A4F498E",
            INIT_RAM_1B => X"EF352A083BBC14A02088E2080C0E0264924902A0029B50370AA40BA33F631ACF",
            INIT_RAM_1C => X"452F48BD26CC14BD22F49B3352B48BD263052B48BD26D2E8BACDF3782E24A80E",
            INIT_RAM_1D => X"04112CC112E82E81E2CCD48D22F498E92EEF052DB3BBC14AD4CC14AD22F49B30",
            INIT_RAM_1E => X"00E229D210C1DD0DC1DD0EC1DD0EC1DD3CF07743E52802B084A003A01BC7CB4B",
            INIT_RAM_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01",
            INIT_RAM_20 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555555555555555555555555555555",
            INIT_RAM_21 => X"AAAAAAAAFFFFFFFFAAAAAAAAAAAAAAAA55555555555555550000000000000000",
            INIT_RAM_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_24 => X"AAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAA5555555555555555",
            INIT_RAM_25 => X"AAAAAAAAFFFFFFFFFFFFFFFF55555555FFFFFFFFFFFFFFFFFFFFFFFF55555555",
            INIT_RAM_26 => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_27 => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_2B => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050",
            INIT_RAM_2F => X"FEFEFAFA54545050FEFEFAFAFEFEFAFAFEFEFAFA54545050FEFEFAFAFEFEFAFA",
            INIT_RAM_30 => X"555500000000FFFF555500000000FFFFFFFFFFFFFFFFFFFFFFFFEB02567E5018",
            INIT_RAM_31 => X"FFFFAAAA5555FFFFFFFFAAAA5555FFFFFFFFAAAAFFFFFFFFFFFFAAAAFFFFFFFF",
            INIT_RAM_32 => X"E7E7EFEF4143FFFFE7E7EFEF4343FFFFE7E7EFEF4243FFFFE7E7EFEF4343FFFF",
            INIT_RAM_33 => X"E7E7EFEF4243FFFFE7E7EFEF4243FFFFE7E7EFEF4143FFFFE7E7EFEF4143FFFF",
            INIT_RAM_34 => X"000000000000FFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_35 => X"FFFF00000000FFFF000000000000FFFF000000000000FFFF00000000FFFFFFFF",
            INIT_RAM_36 => X"FF5FFF5FFF5FFF5FAA0FAA0FAA0FAA0F5F0F5F0F5F0F5F0FFFFFFFFFFFFFFFFF",
            INIT_RAM_37 => X"FF5FFF5FFF5FFF5FAA0FAA0FAA0FAA0F5F0F5F0F5F0F5F0FFFFFFFFFFFFFFFFF",
            INIT_RAM_38 => X"C303030F0303FFFFC303030F0303FFFFC303030F0303FFFFC303030F0303FFFF",
            INIT_RAM_39 => X"C303030F0303FFFFC303030F0303FFFFC303030F0303FFFFC303030F0303FFFF",
            INIT_RAM_3A => X"C00FC00FC00FC00F000F000F000F000F030F030F030F030FFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFF6555544473322211100005757575746464575646757467467467567567564",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3F => X"03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"ADB65323690E3D62284DD8DC280CE238C8CD8C8E231882961965A65B61861865",
            INIT_RAM_01 => X"4E3888A2A0ADA08A82B66828A22208A04242D288802B5A490A79226820FE2E89",
            INIT_RAM_02 => X"94D222322B62223B6D2392508E26B22288A0839300B1E1A023389CEA2288A22A",
            INIT_RAM_03 => X"8A20AD8A0B602A28A0B602A28A0B422A2882B6222FED822E0B0020BADB73AEB2",
            INIT_RAM_04 => X"8C8A2223B48E4862208E26B222B4A538E588823388B0B6D0AD8220AD80A20AD8",
            INIT_RAM_05 => X"6088C3D80A230F62288C3D88C3834A8A2B0E0D2A28AC30D8A8A2B0F622224A08",
            INIT_RAM_06 => X"8BC5242B5F8CC42B64E6288B00BDF4DCA2281B89289888CE23F630A19622230F",
            INIT_RAM_07 => X"8992B88AEAD2B1188ADA9ECC2B422B10AD8AC42B4A2B10ADF1080AD208A60AD2",
            INIT_RAM_08 => X"888AA083F8A2289AD24A0B000002E48448802270B0222222738AA2227F8AA330",
            INIT_RAM_09 => X"88A02B8AE22222D4E8B48B88AE389222A6E988DDBC2F3CA0AD909E48BAA6A9A0",
            INIT_RAM_0A => X"C8498F2126290CA5226909A42B4ADC888888B223F232A32A32A32284888A8270",
            INIT_RAM_0B => X"32122849888A8280AE2BBE8D4C02D581D60338898CD98232362222FC849B2126",
            INIT_RAM_0C => X"280AE2B88888B53A0FB8B58222B4A2888FB8888888B1223F2321A2321A2321A2",
            INIT_RAM_0D => X"F36290CA12F76909A428612222332CCC8FC8CCE8CCE8CCE8CCCA973222A09C22",
            INIT_RAM_0E => X"EBAC9425A08A4CA648A29A2608A6A622B4823362222FC84CDB21336C87CD8F21",
            INIT_RAM_0F => X"8A2A00008BC0000803188D1A22488444A2348AE63722C88888E32273AEB2509C",
            INIT_RAM_10 => X"0023BF0020B02D5A820082E2F00082CF88200BE3000882C0BD002F7000CD8220",
            INIT_RAM_11 => X"086A03C7C7CEA03EBAA4CFCA2C787EEA0B602C08E2981207F0020802082FC03F",
            INIT_RAM_12 => X"64A81208EE70E4EA7C7A0AAF93E7C4D1EB0E7CF56A038C78D7CC7C7C7A0AAAEA",
            INIT_RAM_13 => X"7A0AA4B7AB079C0CE8FFCE70C79C347EEB930B9C3C6A5F1B0A3C0EAC39CE9F0A",
            INIT_RAM_14 => X"888BC2A06AE23C22338A20A422089DCC8DE93794DCCBFDE223309CC6E706FECC",
            INIT_RAM_15 => X"F02237F8A2233948A22888CC223118DEC8DEC8DD55A2338BCFA2E882338BAAB1",
            INIT_RAM_16 => X"A0AA58B80B9F5F3EADB8862F1AB6AB78CC23708CF81236308CFD9590C8C8FDF1",
            INIT_RAM_17 => X"CE222E7CA0880F00B8FBA0ABAA8A2D48618D2083918AA2E0000022C62AF38822",
            INIT_RAM_18 => X"9B25E8CBD8BC6A2B4AA8EF60B8C8C6A0F2376909A42B8AEF0B622008A2672290",
            INIT_RAM_19 => X"21080822F00A4C2A2108048BC028A689822884202BC02B884200A08B90822198",
            INIT_RAM_1A => X"D28028AD248AB44442B7918B98CC26282AA00A92A62390E7C25F0082029F00A2",
            INIT_RAM_1B => X"208828440C82A0A188A2E88A8A8A2A00000022C62A83CE208B80894A2B4A028A",
            INIT_RAM_1C => X"A82300BC0221A08C02F0088482B00BC028A82B00BC02262A0A2B8AE8A646A103",
            INIT_RAM_1D => X"483AA212AA28AC222A21209C02F00B370320A82700C82A082221A0AC02F00886",
            INIT_RAM_1E => X"62288AE9C8EEAEA8EEAEA8EEAEA8EEAE8A3BABAA2A2A8A8C90A188A132CEE888",
            INIT_RAM_1F => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E",
            INIT_RAM_20 => X"AAAAAAAAAAAAAAAA5555555555555555AAAAAAAAAAAAAAAA5555555555555555",
            INIT_RAM_21 => X"AAAAAAAAFFFFFFFFFFFFFFFF55555555FFFFFFFFFFFFFFFFFFFFFFFF55555555",
            INIT_RAM_22 => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_23 => X"65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE65E5EEEE",
            INIT_RAM_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_26 => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_27 => X"7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A7FAA5F0A",
            INIT_RAM_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2A => X"FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050FEFEFAFA54545050",
            INIT_RAM_2B => X"FEFEFAFA54545050FEFEFAFAFEFEFAFAFEFEFAFA54545050FEFEFAFAFEFEFAFA",
            INIT_RAM_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_2E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55555555555555555555555555555555",
            INIT_RAM_2F => X"AAAAAAAAFFFFFFFFAAAAAAAAAAAAAAAA55555555555555550000000000000000",
            INIT_RAM_30 => X"55555555FFFFFFFF00000000AAAAFFFFFFFFFFFFFFFFFFFFFFFFC05401150004",
            INIT_RAM_31 => X"FFFFFFFFFFFFFFFFAAAAAAAAAAAAFFFF55555555FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_32 => X"FFAB5F0F5D0BFFFFFFAB5F0F5C0BFFFFFFAB5F0F5C0BFFFFFFAB5F0F5C0BFFFF",
            INIT_RAM_33 => X"FFAB5F0F5D0BFFFFFFAB5F0F5C0BFFFFFFAB5F0F5C0BFFFFFFAB5F0F5D0BFFFF",
            INIT_RAM_34 => X"000000000000FFFF000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_35 => X"FFFF00000000FFFF000000000000FFFF000000000000FFFF00000000FFFFFFFF",
            INIT_RAM_36 => X"A00FA00FA00FA00FA00FA00FA00FA00FAFAFAFAFAFAFAFAFFFFFFFFFFFFFFFFF",
            INIT_RAM_37 => X"F55FF55FF55FF55FF55FF55FF55FF55FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_38 => X"C303030F0303FFFFC303030F0303FFFFC303030F0303FFFFC303030F0303FFFF",
            INIT_RAM_39 => X"C303030F0303FFFFC303030F0303FFFFC303030F0303FFFFC303030F0303FFFF",
            INIT_RAM_3A => X"C00FC00FC00FC00F000F000F000F000F030F030F030F030FFFFFFFFFFFFFFFFF",
            INIT_RAM_3B => X"FFF98BA98BA8BA98BA98BA98BAA9988BBAA998BBAA988BBA998BBA998BBA9988",
            INIT_RAM_3C => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3E => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3F => X"03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_3_AD_i
        );

end Behavioral; --Gowin_pROM_1541_8k_rom
