--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Thu Sep 21 21:33:04 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_chargen is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(11 downto 0)
    );
end Gowin_pROM_chargen;

architecture Behavioral of Gowin_pROM_chargen is

    signal prom_inst_0_dout_w: std_logic_vector(27 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(27 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(3 downto 0) <= prom_inst_0_DO_o(3 downto 0) ;
    prom_inst_0_dout_w(27 downto 0) <= prom_inst_0_DO_o(31 downto 4) ;
    prom_inst_1_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(7 downto 4) <= prom_inst_1_DO_o(3 downto 0) ;
    prom_inst_1_dout_w(27 downto 0) <= prom_inst_1_DO_o(31 downto 4) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 4,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0C66E06C0000800E0E00800E08C666C80C60006C0C66C66C0666E6C80C20EE6C",
            INIT_RAM_01 => X"0C66666C066EEE660333BF730E00000006C808C608CCCCCE0C88888C0666E666",
            INIT_RAM_02 => X"037FB33308C666660C6666660888888E0C66C06C06C8C66C0EC6666C0000C66C",
            INIT_RAM_03 => X"000FF0008888EC800CCCCCCC0C20C02C0C00000C0E008C6E0888C666066C8C66",
            INIT_RAM_04 => X"000008C60F678C6C06608C6208C6C0E8066F6F66000006660800888800000000",
            INIT_RAM_05 => X"0008C630088000000000E000088000000088E880006CFC60008CCC800C80008C",
            INIT_RAM_06 => X"08888C6E0C66C06C0C666C0E066F6EE60C66C66C0E00C66C0E8888880C666E6C",
            INIT_RAM_07 => X"0808C66C008C6C80000E0E000E80008E08800800008008000C66E66C0C66C66C",
            INIT_RAM_08 => X"0000000000FF000000000FF00000FF00000FF000888888880ECFFEC8000FF000",
            INIT_RAM_09 => X"000000FF0008CE7337EC8000FF000000000008880007FC8888800000CCCCCCCC",
            INIT_RAM_0A => X"0CE66EC037ECCE7388CF70000000000008CEFFF60FF000000CEEEEC0333333FF",
            INIT_RAM_0B => X"137FFFFF0666E3008888888800000000888FF88808CEFEC8666666660C886688",
            INIT_RAM_0C => X"3333333333CC33CC00000000F00000000000000FFFFF00000000000000000000",
            INIT_RAM_0D => X"FF00000088888000000FF888FFFF0000888FF8883333333300008CEF33CC0000",
            INIT_RAM_0E => X"000000FF77777777000000000000000088888888888FF000000FF888888FF000",
            INIT_RAM_0F => X"FFFF000000000000000888880000FFFF00000000FF333333FFF0000000000FFF",
            INIT_RAM_10 => X"F3991F93FFFF7FF1F1FF7FF1F7399937F39FFF93F3993993F9991937F39F1193",
            INIT_RAM_11 => X"F3999993F9911199FCCC408CF1FFFFFFF937F739F7333331F3777773F9991999",
            INIT_RAM_12 => X"FC804CCCF7399999F3999999F7777771F3993F93F9373993F1399993FFFF3993",
            INIT_RAM_13 => X"FFF00FFF7777137FF3333333F3DF3FD3F3FFFFF3F1FF7391F7773999F9937399",
            INIT_RAM_14 => X"FFFFF739F0987393F99F739DF7393F17F9909099FFFFF999F7FF7777FFFFFFFF",
            INIT_RAM_15 => X"FFF739CFF77FFFFFFFFF1FFFF77FFFFFFF77177FFF93039FFF73337FF37FFF73",
            INIT_RAM_16 => X"F7777391F3993F93F39993F1F9909119F3993993F1FF3993F1777777F3999193",
            INIT_RAM_17 => X"F7F73993FF73937FFFF1F1FFF17FFF71F77FF7FFFF7FF7FFF3991993F3993993",
            INIT_RAM_18 => X"FFFFFFFFFF00FFFFFFFFF00FFFFF00FFFFF00FFF77777777F1300137FFF00FFF",
            INIT_RAM_19 => X"FFFFFF00FFF7318CC8137FFF00FFFFFFFFFFF777FFF80377777FFFFF33333333",
            INIT_RAM_1A => X"F319913FC813318C77308FFFFFFFFFFFF7310009F00FFFFFF311113FCCCCCC00",
            INIT_RAM_1B => X"EC800000F9991CFF77777777FFFFFFFF77700777F731013799999999F3779977",
            INIT_RAM_1C => X"CCCCCCCCCC33CC33FFFFFFFF0FFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_1D => X"00FFFFFF77777FFFFFF007770000FFFF77700777CCCCCCCCFFFF7310CC33FFFF",
            INIT_RAM_1E => X"FFFFFF0088888888FFFFFFFFFFFFFFFF7777777777700FFFFFF0077777700FFF",
            INIT_RAM_1F => X"0000FFFFFFFFFFFFFFF77777FFFF0000FFFFFFFF00CCCCCC000FFFFFFFFFF000",
            INIT_RAM_20 => X"C6E66E000888E8E00C0E6C000E66E6600C000C000C66C0000E6E6C000C20EE6C",
            INIT_RAM_21 => X"0C666C0006666C0003BFF6000C88888006C8C000C66660600C8880800666C000",
            INIT_RAM_22 => X"06EFB30008C666000E6666000E888E800C6C0E0000006C0066E66E0000C66C00",
            INIT_RAM_23 => X"000FF0008888EC800CCCCCCC0C20C02C0C00000C0E08CE008CE6660006C8C600",
            INIT_RAM_24 => X"000008C60F678C6C06608C6208C6C0E8066F6F66000006660800888800000000",
            INIT_RAM_25 => X"0008C630088000000000E000088000000088E880006CFC60008CCC800C80008C",
            INIT_RAM_26 => X"08888C6E0C66C06C0C666C0E066F6EE60C66C66C0E00C66C0E8888880C666E6C",
            INIT_RAM_27 => X"0808C66C008C6C80000E0E000E80008E08800800008008000C66E66C0C66C66C",
            INIT_RAM_28 => X"0C66E06C0000800E0E00800E08C666C80C60006C0C66C66C0666E6C8000FF000",
            INIT_RAM_29 => X"0C66666C066EEE660333BF730E00000006C808C608CCCCCE0C88888C0666E666",
            INIT_RAM_2A => X"037FB33308C666660C6666660888888E0C66C06C06C8C66C0EC6666C0000C66C",
            INIT_RAM_2B => X"6C936C93CC33CC338888888800000000888FF8880E008C6E0888C666066C8C66",
            INIT_RAM_2C => X"3333333333CC33CC00000000F00000000000000FFFFF00000000000000000000",
            INIT_RAM_2D => X"FF00000088888000000FF888FFFF0000888FF88833333333639C639C33CC0000",
            INIT_RAM_2E => X"000000FF77777777000000000000000088888888888FF000000FF888888FF000",
            INIT_RAM_2F => X"FFFF000000000000000888880000FFFF000000000008C631FFF0000000000FFF",
            INIT_RAM_30 => X"391991FFF777171FF3F193FFF199199FF3FFF3FFF3993FFFF19193FFF39F1193",
            INIT_RAM_31 => X"F39993FFF99993FFFC4009FFF377777FF9373FFF39999F9FF3777F7FF9993FFF",
            INIT_RAM_32 => X"F9104CFFF73999FFF19999FFF177717FF393F1FFFFFF93FF991991FFFF3993FF",
            INIT_RAM_33 => X"FFF00FFF7777137FF3333333F3DF3FD3F3FFFFF3F1F731FF731999FFF93739FF",
            INIT_RAM_34 => X"FFFFF739F0987393F99F739DF7393F17F9909099FFFFF999F7FF7777FFFFFFFF",
            INIT_RAM_35 => X"FFF739CFF77FFFFFFFFF1FFFF77FFFFFFF77177FFF93039FFF73337FF37FFF73",
            INIT_RAM_36 => X"F7777391F3993F93F39993F1F9909119F3993993F1FF3993F1777777F3999193",
            INIT_RAM_37 => X"F7F73993FF73937FFFF1F1FFF17FFF71F77FF7FFFF7FF7FFF3991993F3993993",
            INIT_RAM_38 => X"F3991F93FFFF7FF1F1FF7FF1F7399937F39FFF93F3993993F9991937FFF00FFF",
            INIT_RAM_39 => X"F3999993F9911199FCCC408CF1FFFFFFF937F739F7333331F3777773F9991999",
            INIT_RAM_3A => X"FC804CCCF7399999F3999999F7777771F3993F93F9373993F1399993FFFF3993",
            INIT_RAM_3B => X"936C936C33CC33CC77777777FFFFFFFF77700777F1FF7391F7773999F9937399",
            INIT_RAM_3C => X"CCCCCCCCCC33CC33FFFFFFFF0FFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"00FFFFFF77777FFFFFF007770000FFFF77700777CCCCCCCC9C639C63CC33FFFF",
            INIT_RAM_3E => X"FFFFFF0088888888FFFFFFFFFFFFFFFF7777777777700FFFFFF0077777700FFF",
            INIT_RAM_3F => X"0000FFFFFFFFFFFFFFF77777FFFF0000FFFFFFFFFFF739CE000FFFFFFFFFF000"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 4,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0366666306667667076676670766666703666663076676670666763103666663",
            INIT_RAM_01 => X"0366666306667776066667760766666606677766036000010311111306667666",
            INIT_RAM_02 => X"0677666601366666036666660111111703603663066776670036666306667667",
            INIT_RAM_03 => X"0137731011117310030000030F63731003333333076310070111366606631366",
            INIT_RAM_04 => X"00000100036633630463106601703631066F6F66000006660100111100000000",
            INIT_RAM_05 => X"06310000011000000000700031100000001171100063F3600310001300133310",
            INIT_RAM_06 => X"0111106703667663036007670007610003601063076300630711131103667663",
            INIT_RAM_07 => X"0101006307100017000707000013631031100100001001000360366303663663",
            INIT_RAM_08 => X"3333333300FF000000000FF00000FF00000FF0001111111103177310000FF000",
            INIT_RAM_09 => X"CCCCCCFFCE731000000137ECFFCCCCCC000EF31100000111113FE00000000000",
            INIT_RAM_0A => X"03766730CE7337EC1110000066666666001377730FF0000003777730000000FF",
            INIT_RAM_0B => X"0000137F033730001111111133CC33CC111FF111001373100000000003116611",
            INIT_RAM_0C => X"0000000033CC33CCCCCCCCCCF00000000000000FFFFF0000FFFFFFFF00000000",
            INIT_RAM_0D => X"FF000000111FF000000111110000000011111111000000008CEFFFFF33CC0000",
            INIT_RAM_0E => X"000000FF00000000EEEEEEEECCCCCCCC111FF111111FF000000FF11111111000",
            INIT_RAM_0F => X"0000FFFF0000FFFF000FF11100000000FFFF0000FF000000FFF0000000000FFF",
            INIT_RAM_10 => X"FC99999CF9998998F8998998F8999998FC99999CF8998998F99989CEFC99999C",
            INIT_RAM_11 => X"FC99999CF9998889F9999889F8999999F9988899FC9FFFFEFCEEEEECF9998999",
            INIT_RAM_12 => X"F9889999FEC99999FC999999FEEEEEE8FC9FC99CF9988998FFC9999CF9998998",
            INIT_RAM_13 => X"FEC88CEFEEEE8CEFFCFFFFFCF09C8CEFFCCCCCCCF89CEFF8FEEEC999F99CEC99",
            INIT_RAM_14 => X"FFFFFEFFFC99CC9CFB9CEF99FE8FC9CEF9909099FFFFF999FEFFEEEEFFFFFFFF",
            INIT_RAM_15 => X"F9CEFFFFFEEFFFFFFFFF8FFFCEEFFFFFFFEE8EEFFF9C0C9FFCEFFFECFFECCCEF",
            INIT_RAM_16 => X"FEEEEF98FC99899CFC9FF898FFF89EFFFC9FEF9CF89CFF9CF8EEECEEFC99899C",
            INIT_RAM_17 => X"FEFEFF9CF8EFFFE8FFF8F8FFFFEC9CEFCEEFFEFFFFEFFEFFFC9FC99CFC99C99C",
            INIT_RAM_18 => X"CCCCCCCCFF00FFFFFFFFF00FFFFF00FFFFF00FFFEEEEEEEEFCE88CEFFFF00FFF",
            INIT_RAM_19 => X"33333300318CEFFFFFFEC81300333333FFF10CEEFFFFFEEEEEC01FFFFFFFFFFF",
            INIT_RAM_1A => X"FC8998CF318CC813EEEFFFFF99999999FFEC888CF00FFFFFFC8888CFFFFFFF00",
            INIT_RAM_1B => X"FFFFEC80FCC8CFFFEEEEEEEECC33CC33EEE00EEEFFEC8CEFFFFFFFFFFCEE99EE",
            INIT_RAM_1C => X"FFFFFFFFCC33CC33333333330FFFFFFFFFFFFFF00000FFFF00000000FFFFFFFF",
            INIT_RAM_1D => X"00FFFFFFEEE00FFFFFFEEEEEFFFFFFFFEEEEEEEEFFFFFFFF73100000CC33FFFF",
            INIT_RAM_1E => X"FFFFFF00FFFFFFFF1111111133333333EEE00EEEEEE00FFFFFF00EEEEEEEEFFF",
            INIT_RAM_1F => X"FFFF0000FFFF0000FFF00EEEFFFFFFFF0000FFFF00FFFFFF000FFFFFFFFFF000",
            INIT_RAM_20 => X"7036630001113100036763000366300003666300076676600363030003666663",
            INIT_RAM_21 => X"0366630006666700066776000311113006676660300000000311301006667660",
            INIT_RAM_22 => X"0337660001366600036666000011171007036300066667000036630066766700",
            INIT_RAM_23 => X"0137731011117310030000030F63731003333333073107007036660006313600",
            INIT_RAM_24 => X"00000100036633630463106601703631066F6F66000006660100111100000000",
            INIT_RAM_25 => X"06310000011000000000700031100000001171100063F3600310001300133310",
            INIT_RAM_26 => X"0111106703667663036007670007610003601063076300630711131103667663",
            INIT_RAM_27 => X"0101006307100017000707000013631031100100001001000360366303663663",
            INIT_RAM_28 => X"03666663066676670766766707666667036666630766766706667631000FF000",
            INIT_RAM_29 => X"0366666306667776066667760766666606677766036000010311111306667666",
            INIT_RAM_2A => X"0677666601366666036666660111111703603663066776670036666306667667",
            INIT_RAM_2B => X"6C936C93CC33CC331111111133CC33CC111FF111076310070111366606631366",
            INIT_RAM_2C => X"0000000033CC33CCCCCCCCCCF00000000000000FFFFF0000FFFFFFFF00000000",
            INIT_RAM_2D => X"FF000000111FF00000011111000000001111111100000000639C639C33CC0000",
            INIT_RAM_2E => X"000000FF00000000EEEEEEEECCCCCCCC111FF111111FF000000FF11111111000",
            INIT_RAM_2F => X"0000FFFF0000FFFF000FF11100000000FFFF000006776000FFF0000000000FFF",
            INIT_RAM_30 => X"8FC99CFFFEEECEFFFC989CFFFC99CFFFFC999CFFF899899FFC9CFCFFFC99999C",
            INIT_RAM_31 => X"FC999CFFF99998FFF99889FFFCEEEECFF998999FCFFFFFFFFCEECFEFF999899F",
            INIT_RAM_32 => X"FCC899FFFEC999FFFC9999FFFFEEE8EFF8FC9CFFF99998FFFFC99CFF998998FF",
            INIT_RAM_33 => X"FEC88CEFEEEE8CEFFCFFFFFCF09C8CEFFCCCCCCCF8CEF8FF8FC999FFF9CEC9FF",
            INIT_RAM_34 => X"FFFFFEFFFC99CC9CFB9CEF99FE8FC9CEF9909099FFFFF999FEFFEEEEFFFFFFFF",
            INIT_RAM_35 => X"F9CEFFFFFEEFFFFFFFFF8FFFCEEFFFFFFFEE8EEFFF9C0C9FFCEFFFECFFECCCEF",
            INIT_RAM_36 => X"FEEEEF98FC99899CFC9FF898FFF89EFFFC9FEF9CF89CFF9CF8EEECEEFC99899C",
            INIT_RAM_37 => X"FEFEFF9CF8EFFFE8FFF8F8FFFFEC9CEFCEEFFEFFFFEFFEFFFC9FC99CFC99C99C",
            INIT_RAM_38 => X"FC99999CF9998998F8998998F8999998FC99999CF8998998F99989CEFFF00FFF",
            INIT_RAM_39 => X"FC99999CF9998889F9999889F8999999F9988899FC9FFFFEFCEEEEECF9998999",
            INIT_RAM_3A => X"F9889999FEC99999FC999999FEEEEEE8FC9FC99CF9988998FFC9999CF9998998",
            INIT_RAM_3B => X"936C936C33CC33CCEEEEEEEECC33CC33EEE00EEEF89CEFF8FEEEC999F99CEC99",
            INIT_RAM_3C => X"FFFFFFFFCC33CC33333333330FFFFFFFFFFFFFF00000FFFF00000000FFFFFFFF",
            INIT_RAM_3D => X"00FFFFFFEEE00FFFFFFEEEEEFFFFFFFFEEEEEEEEFFFFFFFF9C639C63CC33FFFF",
            INIT_RAM_3E => X"FFFFFF00FFFFFFFF1111111133333333EEE00EEEEEE00FFFFFF00EEEEEEEEFFF",
            INIT_RAM_3F => X"FFFF0000FFFF0000FFF00EEEFFFFFFFF0000FFFFF9889FFF000FFFFFFFFFF000"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

end Behavioral; --Gowin_pROM_chargen
