--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.9.02
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Thu Apr 25 13:22:34 2024

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_SDPB_kernal_8k is
    port (
        dout: out std_logic_vector(7 downto 0);
        clka: in std_logic;
        cea: in std_logic;
        reseta: in std_logic;
        clkb: in std_logic;
        ceb: in std_logic;
        resetb: in std_logic;
        oce: in std_logic;
        ada: in std_logic_vector(12 downto 0);
        din: in std_logic_vector(7 downto 0);
        adb: in std_logic_vector(12 downto 0)
    );
end Gowin_SDPB_kernal_8k;

architecture Behavioral of Gowin_SDPB_kernal_8k is

    signal sdpb_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal sdpb_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal sdpb_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal sdpb_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal sdpb_inst_0_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_0_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_0_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_0_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_0_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_1_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_1_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_1_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_1_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_1_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_2_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_2_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_2_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_2_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_2_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_3_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_3_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_3_ADA_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_3_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_3_ADB_i: std_logic_vector(13 downto 0);
    signal sdpb_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component SDPB
        generic (
            READ_MODE: in bit := '0';
            BIT_WIDTH_0: in integer :=16;
            BIT_WIDTH_1: in integer :=16;
            BLK_SEL_0: in bit_vector := "000";
            BLK_SEL_1: in bit_vector := "000";
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLKA: in std_logic;
            CEA: in std_logic;
            RESETA: in std_logic;
            CLKB: in std_logic;
            CEB: in std_logic;
            RESETB: in std_logic;
            OCE: in std_logic;
            BLKSELA: in std_logic_vector(2 downto 0);
            BLKSELB: in std_logic_vector(2 downto 0);
            ADA: in std_logic_vector(13 downto 0);
            DI: in std_logic_vector(31 downto 0);
            ADB: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    sdpb_inst_0_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_0_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_0_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_0_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(1 downto 0);
    sdpb_inst_0_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= sdpb_inst_0_DO_o(1 downto 0) ;
    sdpb_inst_0_dout_w(29 downto 0) <= sdpb_inst_0_DO_o(31 downto 2) ;
    sdpb_inst_1_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_1_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_1_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_1_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(3 downto 2);
    sdpb_inst_1_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= sdpb_inst_1_DO_o(1 downto 0) ;
    sdpb_inst_1_dout_w(29 downto 0) <= sdpb_inst_1_DO_o(31 downto 2) ;
    sdpb_inst_2_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_2_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_2_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_2_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(5 downto 4);
    sdpb_inst_2_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= sdpb_inst_2_DO_o(1 downto 0) ;
    sdpb_inst_2_dout_w(29 downto 0) <= sdpb_inst_2_DO_o(31 downto 2) ;
    sdpb_inst_3_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_3_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_3_ADA_i <= ada(12 downto 0) & gw_gnd;
    sdpb_inst_3_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(7 downto 6);
    sdpb_inst_3_ADB_i <= adb(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= sdpb_inst_3_DO_o(1 downto 0) ;
    sdpb_inst_3_dout_w(29 downto 0) <= sdpb_inst_3_DO_o(31 downto 2) ;

    sdpb_inst_0: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"1445216085A804D5F21600D120DE21490D113070306524545614C534083054C9",
            INIT_RAM_01 => X"CA8B00E31445644B47A9658C09801780D3164D901926432BC0C30902100E0132",
            INIT_RAM_02 => X"2C9CD03A5091144C361903D38DB10038DB13D245F28030238004D3C038E09210",
            INIT_RAM_03 => X"E18A063860818B28510B41133C590CC24B1CA18E32662274C64DF0E30726707C",
            INIT_RAM_04 => X"44003CA8500C81D32AC628A385A2828E04C50A828530A6E24D070C1240204E28",
            INIT_RAM_05 => X"D473CB68403ADEB590F0260991E03480AB247832370C0C89C276524442408933",
            INIT_RAM_06 => X"1C001EAF4292A0D9B4017E2F003D89DFB30C0081C50CC9F107145C309ADCD677",
            INIT_RAM_07 => X"649661D11DD0B7920D4985C5E3581C444BC041306261E8A0B88F0C030CB0228D",
            INIT_RAM_08 => X"F2A801C568D18DD8CCB137AB390FE0E005411B4DE03400D0A3B400E0ED00EC0A",
            INIT_RAM_09 => X"111475155531404936931761A04562022B7B490B4100A3C90305AA28DD821B35",
            INIT_RAM_0A => X"500B4404DA8C089C25DC80411210611519669986D1876D1D94503290CAC10802",
            INIT_RAM_0B => X"5CCA926860D72CC0BA434CA467800A482D84AC32F41E519D610014D205804843",
            INIT_RAM_0C => X"89D08D5E332A319447020E1802018CEDD5CC120C81D98442B143280030C15040",
            INIT_RAM_0D => X"D102904B15445945466AA23129CCA6373578C0080281A2CA8A0863849151090D",
            INIT_RAM_0E => X"24DA54710D3451483013CD2081B30AC8363404044C5C3370440B43110A903A28",
            INIT_RAM_0F => X"CCC0154C1C213164C198DD80CA000D01A805A041168C002910C30C56337626CC",
            INIT_RAM_10 => X"A630C1A108DA34A3011085D1094423404DACA85B050A82DA54730D3451481140",
            INIT_RAM_11 => X"1D6AE349141E4E5B8C42A020278A84A22133768A2213346A8038B8890A052310",
            INIT_RAM_12 => X"8AA6202026C528114934AA515515C014623549C0424450040D9670445C101114",
            INIT_RAM_13 => X"098755413475646010D951C4161D4289829184D9C939C44044D0891098D24506",
            INIT_RAM_14 => X"5B17560405402056019AADD827916EEC514641E011D9D5365C20592205122043",
            INIT_RAM_15 => X"3535228D8E07125CB00060CB1032259434154880514206675544C181C0944200",
            INIT_RAM_16 => X"0FB609E575A606E01905258A536501DA2D892A84A244C022C08BB22481041414",
            INIT_RAM_17 => X"88DE5D12E43BD2592370B895E1F7914F623797E0290EF49648DC2E25787DE450",
            INIT_RAM_18 => X"FFFBA2597615251C1A0150725241C9FE137977038BA5C660F79F12167392353D",
            INIT_RAM_19 => X"0000000077D739390E68003000F000000003DF78EF94CFC3BDA692B70B88DEDC",
            INIT_RAM_1A => X"92CC811B2045151A324C93248C902440B2CA044516305814E243880041040000",
            INIT_RAM_1B => X"D35114680144042100324918E01144751116020D0402489145354D10644751AA",
            INIT_RAM_1C => X"A30200648114492045151868064818945009324516C354D5C924512C924AA614",
            INIT_RAM_1D => X"210941DD9700723173CF0C4008CC1D00860922881144445111D44445111D4401",
            INIT_RAM_1E => X"80A004150047853000E2008520B022B25585210A8E21382A5585210834011485",
            INIT_RAM_1F => X"200C5210BCF1693C482152C521085053568C211A0856C8D511531845013CA0C8",
            INIT_RAM_20 => X"27370507C0621464C03406A0B72A4149F282BB8DE0727DC9E72546E929460020",
            INIT_RAM_21 => X"503618510404350B6D412E3939772E93D734DD100E1C218C030A61B6C1574716",
            INIT_RAM_22 => X"5068F0281514DA16677140010444089050C0E341511F4279E5999399DE471D24",
            INIT_RAM_23 => X"F08527150427C500BC1403803642555DDA5DB01406432500003C002005E01850",
            INIT_RAM_24 => X"150888D0C00944DD327CD33CF20272042154A9348FE181433627CD33CD208644",
            INIT_RAM_25 => X"594000A284316A8204411C1224062D1D03478010EC13303424BC08C3C8094C61",
            INIT_RAM_26 => X"12362D995456512B320A8CF38C21469CC463238445966D194095228442596DB6",
            INIT_RAM_27 => X"4D00DF01054154244632142180C701310C4878031010C8A7170585B10714FCCD",
            INIT_RAM_28 => X"8C1C00047418888C1D7050620619DD4CB81122C2E00AA5E1C6995DCB815A08C1",
            INIT_RAM_29 => X"CCD0456CD19D0B6C0A19B1C55274517184CC44DF32447700E891C84E1C130D88",
            INIT_RAM_2A => X"82D0001534E10348B36D188428080923045344304A1CC0E8A92010900C8286B2",
            INIT_RAM_2B => X"C55C4DF32789551B29C48D4230E34031CC4D70214CA016F1C860118DD022E2A8",
            INIT_RAM_2C => X"509111084B66A080914818507550944610C01A33450604F1541E0145426CD30C",
            INIT_RAM_2D => X"914270335401A406905801010609B20145A628D195590A1A2894713143C04153",
            INIT_RAM_2E => X"84415207B000201610E251CC500C5C118152C067480381072103014134914134",
            INIT_RAM_2F => X"71C91D5997344130B73414124CC3124411440CC1C9933408CDB0219410184EC4",
            INIT_RAM_30 => X"4564242041AC8060091064751C4180011108048417200801CC82050E140215C8",
            INIT_RAM_31 => X"51489416601106080000C834026D058C48E4E0D03898913432A880DAA0401624",
            INIT_RAM_32 => X"1D84501605657690641220040658510926055354DD0255C9050CD8DD06402024",
            INIT_RAM_33 => X"B065A914881D94504C5040760DAB170661861018100B511A59B1100911AC4131",
            INIT_RAM_34 => X"F38C45340D4367557602C048D2A15433924245E01C9880025BCA8026D5E358AA",
            INIT_RAM_35 => X"C9B8459D6744D18AD6744D12758954B40A291A714201021460CDC60347262041",
            INIT_RAM_36 => X"D08014181846D5D63904C9450607446150762417021640F6320112128060A84C",
            INIT_RAM_37 => X"089C1527446072038B1CD526805E28010877270741334E141E2A01559820828D",
            INIT_RAM_38 => X"CD5016340041D1C5843057C6207203E96C0D348D334528020B38192CAC8B06CA",
            INIT_RAM_39 => X"0F1441C280CA08E1A08D591051510019B57176007080505D205114200472062E",
            INIT_RAM_3A => X"05D15756484132B08086124151AF6967F8A9EBA910C7714DC0E1081B12C35D60",
            INIT_RAM_3B => X"03B7816415704158A475759D474A8278E274D64910551764C4211A4642202A40",
            INIT_RAM_3C => X"462415C2107140A2023180515D02300A26A26820BA0BA09411150B44B52644A1",
            INIT_RAM_3D => X"8BB3083D082D84103850B4C6541E274080565000849E4C84088241C4A332A28B",
            INIT_RAM_3E => X"A09512455529517094301305180821045050A5508B31BA81E072E00E06EC550C",
            INIT_RAM_3F => X"C2B6A41852CC38C24814238C38C38C38520B14418714B24B2091C52061441CF3"
        )
        port map (
            DO => sdpb_inst_0_DO_o,
            CLKA => clka,
            CEA => cea,
            RESETA => reseta,
            CLKB => clkb,
            CEB => ceb,
            RESETB => resetb,
            OCE => oce,
            BLKSELA => sdpb_inst_0_BLKSELA_i,
            BLKSELB => sdpb_inst_0_BLKSELB_i,
            ADA => sdpb_inst_0_ADA_i,
            DI => sdpb_inst_0_DI_i,
            ADB => sdpb_inst_0_ADB_i
        );

    sdpb_inst_1: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"460684681110A1509046B063286A044A2D2231B480552911948A0297C90287C5",
            INIT_RAM_01 => X"7C0A7089048454945445456402A03A00A0D4210850841047004E04A258450E90",
            INIT_RAM_02 => X"C494D3664492C84E2B7440F8F3CF878F3CF8F9A250F03413431C5FC230EE8079",
            INIT_RAM_03 => X"EE680238900081040023C22C309208C085D071BB01B7F0A57C4ED0BC190A50B4",
            INIT_RAM_04 => X"4BCF24D06F2402FC450F0C13899A004E20090900403229700F0BB423C28087CC",
            INIT_RAM_05 => X"4A9A66E54032E0B83EBC38C152801840C204A80C3B40A40AD0786168C9600A83",
            INIT_RAM_06 => X"2F0002AD3FA4F8389F1723E7F0C95E306370A00242800EB2390A1D0252E27534",
            INIT_RAM_07 => X"83CF09192128843C510A55020C30A0D7A1C0A2B0A2A39094A103105DF0830981",
            INIT_RAM_08 => X"C2A8030D4416020044835E3559D097B10BCD9A65B1098D93426205195E2D9F25",
            INIT_RAM_09 => X"336CEB3FF3105212007FC590620C6AA0B1C1882B8800C0DE8F4FAA042005137F",
            INIT_RAM_0A => X"A0486A89155108AC89E08A0AA6288BDDE2E87E2CB60E8FAD0C90055C154220C0",
            INIT_RAM_0B => X"EC487DD6802420D01F73640F5542A545872C0712FFBC92925D09C3AE754AA499",
            INIT_RAM_0C => X"0E5AA5E500250278492541204542055E50101AA8891909F16254430992020158",
            INIT_RAM_0D => X"12B16388256A5A4A69955A1216700C3B054602AAA9095201D42481482525822E",
            INIT_RAM_0E => X"5C01C0B16082082906813412C65C25353839080A30E5C1444AA96055C5B28514",
            INIT_RAM_0F => X"C41420546C58C39302E0EEBE87EC814A58C55AAB09F10B16161824E500940970",
            INIT_RAM_10 => X"59FE827D4427D07C68220E5242472052A1545425C925F901C0B0608208291644",
            INIT_RAM_11 => X"3E95CB6DB6DAA54FFF407224AF0508512A90580512A90481FB055641F549A022",
            INIT_RAM_12 => X"B587A332078994DB6DB655929121C8A4827A42CCA2773C882CBD519B306466CF",
            INIT_RAM_13 => X"012CA473368B7764120C0C4834B2AD81F29209E9C1D2C8A277FCC1E0A2DB6DB5",
            INIT_RAM_14 => X"F907850608442086C2D1C709374007D1D64D8DE05A21110201A4D2A120262481",
            INIT_RAM_15 => X"3A3A10BE480916493ECCEACA02A40F3E0B1924A33CE8CF9694A0CCF3903C8AAB",
            INIT_RAM_16 => X"B22235AD6B982A9CB22F03C3D08F33E58742D6CC3CF59C94B442E0F43D093A19",
            INIT_RAM_17 => X"01CFC32EBF2FB2A5899945112442AFDC0073F0AF2FCBECA962665144491056F7",
            INIT_RAM_18 => X"FFFF7C30FB2A0324A7CBE2E3A08B4EC8173F0FB6F76844B9E5B2EC83D0443F30",
            INIT_RAM_19 => X"88888888C833D540101C0034806000000003CF74FF3FCBF3FB2858DB94D3D2C7",
            INIT_RAM_1A => X"D340C11728CF35AF2388E23881D1388EC34F2CEB3AC1A09615C06859B2C88888",
            INIT_RAM_1B => X"EFB3ACFC896C245914A38D3C62B14CDB3B162BC2C893882FFFFEB7645CCBB3AA",
            INIT_RAM_1C => X"D0070454A33CD528CF35A85F0B4C3324584E10BFFF4FEB728E3458F7D2CA2F30",
            INIT_RAM_1D => X"E33905D1D320322363C70808FD306808040B248A33CCCCB333ECCCCB333ECCA5",
            INIT_RAM_1E => X"4FD7041F104946D010F0228FE0D32343334FC33975007737334FC3380400734F",
            INIT_RAM_1F => X"A220FE2FFFE33D384DAC41FA133CFCA3757C10742B3300DDD241370CF63CF088",
            INIT_RAM_20 => X"28190A0BCC9324A402BE8EA81C2C428EF30A3F0E1CA387461E0B48FA22E4AAAA",
            INIT_RAM_21 => X"290410FC821D38C44E330D1E804C0C13EF20CC3000008200000DC68F8267AA09",
            INIT_RAM_22 => X"F2944E13951824E564624AE93885E454920AC3A3B37BC7777A6171E43793FFCB",
            INIT_RAM_23 => X"F20B0B39080BC00213BF91790A607CF3E1F3CCB904BED4000010012A88B03FF2",
            INIT_RAM_24 => X"27C84A4800290827C24C4C0C5D06D0BF1278AB1071AB0A520924C4C0CFC029C8",
            INIT_RAM_25 => X"B2A5266900F16A960941448D28D55951414B092A542A1308268C2011781B80F1",
            INIT_RAM_26 => X"110A0393E4A4B996C225F031B0924A7C09F02424893E4392C82D298488F38308",
            INIT_RAM_27 => X"C80C55E907829F24491624933B53F3E338B9C9D33834081033CD4D03183B13C1",
            INIT_RAM_28 => X"C70C0D0874A798C491322CB0C4925A40B022A8B8B242CBB044929A4B03D1745B",
            INIT_RAM_29 => X"30C047BBD5D18B700A1DC349E24492724405C824C2448435189A48790C1F8698",
            INIT_RAM_2A => X"8878013812522128B147942CB88A3FCA2560A517843C81D0DCFC28C0C1A286C1",
            INIT_RAM_2B => X"592C824C2431111B74B8018116C20314C44533334DD933E0BDD45D8192955058",
            INIT_RAM_2C => X"BC9122E3E2CF3CC89A48BCE0BA7C909F138224130F3130FF7CDB0389F25C1130",
            INIT_RAM_2D => X"2C897C93848446111810B38CF3CF028CF31114E1A121840504133023497A41E3",
            INIT_RAM_2E => X"0C93A33CC3F2A40512C010C0AE00D4A542CF42654C2B02A32343CABADB6DB6CB",
            INIT_RAM_2F => X"10BD21D214224E6D443421009700218B010100C242891A9B0ABE83242820EC0D",
            INIT_RAM_30 => X"CB3ACA28CD34F0B08B334CFB38CD53FB022C210123E22C80C88B0FEC3A4594C8",
            INIT_RAM_31 => X"FF30BF285022AD2CFCAB04B026227A1951512525B360A2BA82AAA8DDDC8A555C",
            INIT_RAM_32 => X"3E8CE3F52CC7CC7FCBF903F0FCBFA037DF0BFFEB7E71BF42FC80286E2523FBF4",
            INIT_RAM_33 => X"808BA608C4912CB708FC9C2E03A2160ACE05229633C8B32CCD633C8933C8CC07",
            INIT_RAM_34 => X"5D70458A0608494A54C8707CC24266B150B888B0042E22926648080B52C2949A",
            INIT_RAM_35 => X"8A7049951D66B9C951D66B9A7A524A5777CB22E0B0116600A40A06204A08244E",
            INIT_RAM_36 => X"5A48BC202099E94FF1334BCE08CD4A4BE09808BF0A8A8A8B331314F28B3CE888",
            INIT_RAM_37 => X"D2B42E244991FD070C34EE254092144621FA2A0A03160CFB2CEC0D1D1FFC4985",
            INIT_RAM_38 => X"4E5C3A3A3042EA824001557E11B43A66534C2048338650414C302830B04A0700",
            INIT_RAM_39 => X"EE34C301C30C2AC3434DDDD81211E4299652212A30C2F3FEE0320E8B15528550",
            INIT_RAM_3A => X"20E8038040BF8443123820A275D3372100302DD802180640C51B00B01200FF40",
            INIT_RAM_3B => X"3657FDCB76CCB7681C785B3ECDB39BCF30FFFFFFACFFFF9F890B60EBC86A21CA",
            INIT_RAM_3C => X"0CF0CF00D8C340F1C0C300FFFEAA8B80C30C34070C70D01C111D21CA1F0A4999",
            INIT_RAM_3D => X"40D30882C88240A0A7023C8C206CFA02AAFC30B8A534CC8F48AA6300AFC2820B",
            INIT_RAM_3E => X"FFF22FFF2FC722E036073C087AAA1334FC931D7447C30E0951A03805D830C021",
            INIT_RAM_3F => X"ECC804DB5DB3CB2DF5DF7C71C30CF3CBEF3DFBFFFFFFCF39F7DF7EFBEF7CF3EC"
        )
        port map (
            DO => sdpb_inst_1_DO_o,
            CLKA => clka,
            CEA => cea,
            RESETA => reseta,
            CLKB => clkb,
            CEB => ceb,
            RESETB => resetb,
            OCE => oce,
            BLKSELA => sdpb_inst_1_BLKSELA_i,
            BLKSELB => sdpb_inst_1_BLKSELB_i,
            ADA => sdpb_inst_1_ADA_i,
            DI => sdpb_inst_1_DI_i,
            ADB => sdpb_inst_1_ADB_i
        );

    sdpb_inst_2: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"30127BBAECE14E8FCB338269BA6CB32FA829B8BEDB1B499BB20BF24B2D842B24",
            INIT_RAM_01 => X"C61B422DA0B2A0A22AA22ABAA6EA8BA22A22C8B28B22CA23E9FE83A3369826EB",
            INIT_RAM_02 => X"6727DAA8A6028A7DAAAA6808000006820820208AFBC9FA9F29EAF32AF6F28C62",
            INIT_RAM_03 => X"F0A22CBE028B29A2888BE2B07229A3CA6B2E8A89ABAC043AC63EFA92A8C395BE",
            INIT_RAM_04 => X"0B2CB2AAACBAAAF2ABA9A28BE2288A2F8122208A288880DA6F8A0D3AEA84ED22",
            INIT_RAM_05 => X"024F21980039024090C08A6682E89AE22A90B282ABE1BAAAF9318EB212B6AADA",
            INIT_RAM_06 => X"2C8006AC43D1F3BDBCE705C937CFB773CBC1B6AA10A2AECBB840AF84A902989E",
            INIT_RAM_07 => X"630C2448242D36B600EA00E6104E21109409BEEE0F2AE1E97AABA6B3430226E4",
            INIT_RAM_08 => X"0AAAA840124520427D018CA2A6E2209AAB2AEABE9ABA2AAA86A52CCCCDB88DB4",
            INIT_RAM_09 => X"9004392490B60462B42E03B7B60409784138A06B202BB9001020AAB6042F8400",
            INIT_RAM_0A => X"AED1293766442D2E65ED681A56280200200802000212802010AA99AA4439AA62",
            INIT_RAM_0B => X"03D0DAC3250FA602088CBF100A6950D28D3C8EB436FA4242A2AD20E284DA937A",
            INIT_RAM_0C => X"146AA4298C98C989094226031610164E4767601B104252D99C91042034187461",
            INIT_RAM_0D => X"42B92CD0DD296141E5564A859A831BC3D19AE96AA436BA6090D80C82A406189E",
            INIT_RAM_0E => X"61D096A50D3C51CA90AAC8859490DA48B8586162410905990841091AA416905A",
            INIT_RAM_0F => X"0141876D4D6904241861CEE22A2ED41A4B946A9552842B90504B854A85005243",
            INIT_RAM_10 => X"608220A2214A22A10A8D5402149AA506B64F654900DA86D096A50D3C51CA9AAB",
            INIT_RAM_11 => X"0E04E28A28A5554555180B4394A6366B4A4D28A4B4A4D08A8B91010A84D7A85A",
            INIT_RAM_12 => X"440AA84D88D79A8A28A266406C0E969405F9CAEB89E2F36BA0B834292F078A49",
            INIT_RAM_13 => X"A4009D2FA10AA2AAB4DB5BAAA0029262A45017E7129AEB89E2B312AE18A28A2A",
            INIT_RAM_14 => X"2881884860808D8A602080FA809DC206069092EAC426C6B4566A02AB45A9AABA",
            INIT_RAM_15 => X"42F0DC2EDD98C2F20A142B50C0804000C0C3C735048243B2B0ABE49002008AA9",
            INIT_RAM_16 => X"E2228CBF2F8840B14059C6B0140290E08D30883E00202508029024030B60D050",
            INIT_RAM_17 => X"286DC52F74500C25086508605864011C4B1E71E63A18030D431D431C171D0046",
            INIT_RAM_18 => X"FFFCA041BA40C4210A14E584041610C8913715B9DEAEBEBFDB7BDB4E9F500471",
            INIT_RAM_19 => X"72D872D8154800000000000400D000000003DF31D71DC7C7004150455045C545",
            INIT_RAM_1A => X"8A61A8DB4D412828B6AFAB6A1A8AEAF3BA68B4012D0636D2848AB162A88072D8",
            INIT_RAM_1B => X"E99004A2E528816CDA7EA8AEEBD924392D9057628A7EA12492419025841192AA",
            INIT_RAM_1C => X"885AA98F3504AB4D412821AD8A2AAC23A5FA84924A641902DAA28C248AD08BA6",
            INIT_RAM_1D => X"8D2BA0A0AEB6EA85AEAEBA6D4BC18F232DAB4A23504A42129064A411290A4A5A",
            INIT_RAM_1E => X"D4B82369B51BEE324598B6148299E6A652F49D23CFADAA6A52F4BD2258A592F4",
            INIT_RAM_1F => X"8B614A6420F908BED82BEBCDB525499E2BCA8DA94AD01F8A82E8EB642AEA8BA6",
            INIT_RAM_20 => X"73C373E32DCEB1B3A8ECFE0DE6C2F8F8CB252B6E199F06181A59088F42627100",
            INIT_RAM_21 => X"28DBBA4BEFAAB4181D049080041291488390E40AA5825965A4A18042EB328A40",
            INIT_RAM_22 => X"99BED3EC06410B018185AB28E0EB3F2969D8DB8FC58020400104480440000F0A",
            INIT_RAM_23 => X"C804E0C3E1E32888B4A4864841884490E1129248DB8C202222200B436FD8AC99",
            INIT_RAM_24 => X"7A2AD0DFA2945D0C07B6C0F2C1588B0887A2AC9044F4651740FB6C0F2F089C98",
            INIT_RAM_25 => X"51D9D92B2B0D0010D195BAB061A42A42580B6A2621A34CC1F83693DB0562E1B8",
            INIT_RAM_26 => X"85C1C9E272385E6F049BC1CB01E9092A36B8D890AC2F0BC1ED15C610A492C92C",
            INIT_RAM_27 => X"6F23EC285AECE8B90BFBFA61EE000000808F8FBC04084CB108024351ED08741D",
            INIT_RAM_28 => X"6EB6F1D9B6BAEB6306D8288FA2C2CA3D362E84A2DB628ADB22C2CAD36CEB4DC2",
            INIT_RAM_29 => X"C1E91BAC8282122670689A2E8BB6CAEBBE1E5F0D079090E005C253CEB6F36EEB",
            INIT_RAM_2A => X"28DFC8C1FC9B7FC33B06CF1AB2D0FD24518C0BB0DCAA16A1A9B66392362C1A9B",
            INIT_RAM_2B => X"ECA5F0D078E0303A2386362B70DBC8FBA67EE895AAA690FA88810A10AA440209",
            INIT_RAM_2C => X"A2E423A2828A2B65C2526EBA2BA2E7EBA76B2C87A9ADF6A2A6AC8AEE8BB2DB41",
            INIT_RAM_2D => X"28A832071A6223AAAE4190D492439ED41288812A6A2AE86868B0E9B5A70A16BA",
            INIT_RAM_2E => X"04840E8485286AAB50DBCBAAD3616102F24A6B3B36BB6C2E858B20A28A28A28A",
            INIT_RAM_2F => X"EA882A82ABA458B08AF629962C13962C8E698E1038FB62AC308281A10F80EE56",
            INIT_RAM_30 => X"212F0B4148A6D8AAD15224192D4A052D6BFA92126E2B7ADBA67EAC1DBB669BAA",
            INIT_RAM_31 => X"492712668B8EBB8B4AAF617A6833FBB377FB36FB3421CE4AE80036AA90A5AA84",
            INIT_RAM_32 => X"0AF48528A406406409214D2940A8DB50485924190EA992924BED2D029AF92D0F",
            INIT_RAM_33 => X"0606394B670612A05F49AADF7D0859E8B36A296BD230904641B523D0526D4969",
            INIT_RAM_34 => X"92C3149950D10B0B3BA2EBCDEB87394F3443AFD8B2108EDBBB6E3286C6D8AAC0",
            INIT_RAM_35 => X"33363CECDFB33EBECDFB33EF2B0B3B320A0000840FF50996AA50BA990843E210",
            INIT_RAM_36 => X"E598260301ECECFB38D2326226430B02BA08C968A00BD0CC879F8008D92419A1",
            INIT_RAM_37 => X"8A22A8BB6CE4A35B69A2A8BBEFEFBEB89128F073C9FBAD0AAD0CA8282F361E1C",
            INIT_RAM_38 => X"5A4C89527234A2901F3913C88E0000003C1EBA5E8F9B32F679B6ACA6A6D15A62",
            INIT_RAM_39 => X"9DB6DBA5021F97EA86AAAAAE082F362EBBB77CC9DB6AD90EC9445B3091343642",
            INIT_RAM_3A => X"61C0470C2890B30BB4341062EEEEFECDFDCDCCEBB41447136007BBC0B4107328",
            INIT_RAM_3B => X"B333840906F090A32828290E4090144102410410241043A8F280200BA4A64290",
            INIT_RAM_3C => X"AC324BA8A6EB65FBE0872B490E1006E000082180002086024464A1081843ACCC",
            INIT_RAM_3D => X"F1942D0D2D05254F7888BEA2250D2BA2AA40A88D263633B47E6B9BA7AE0EA69B",
            INIT_RAM_3E => X"810424902D0825B56986D0D83C40B52149A802E149031076999C654918605FC6",
            INIT_RAM_3F => X"CEC4582083428A2B4E34D0A28A286186F30C2082CA2493883CE20B34D34D38D0"
        )
        port map (
            DO => sdpb_inst_2_DO_o,
            CLKA => clka,
            CEA => cea,
            RESETA => reseta,
            CLKB => clkb,
            CEB => ceb,
            RESETB => resetb,
            OCE => oce,
            BLKSELA => sdpb_inst_2_BLKSELA_i,
            BLKSELB => sdpb_inst_2_BLKSELB_i,
            ADA => sdpb_inst_2_ADA_i,
            DI => sdpb_inst_2_DI_i,
            ADB => sdpb_inst_2_ADB_i
        );

    sdpb_inst_3: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 2,
            BIT_WIDTH_1 => 2,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"9B2119A06673B666B19A126D206B199A162D2BA8919B3666624CF90ACB0ADA06",
            INIT_RAM_01 => X"123AD2AB1A999899999999A4EA83AA82AF58B62262D8888BC308061149F72691",
            INIT_RAM_02 => X"2326F088BC2209AF088BC424208201020824259EB397BC7BC7B8D7C7BCE58CA6",
            INIT_RAM_03 => X"E5AB0D3862C34D30C08B82F7BC6C12F30960A218298E4CDA1238E18698CD8C38",
            INIT_RAM_04 => X"8AC8206EE824EEE48A8A30C3866AC30E233626C30C08A6A30E0A1F12C54C4A70",
            INIT_RAM_05 => X"89AF080E001B1AC6E5849BC262A09BC26D08ACD7BA8064EEA0B481A405A4EE91",
            INIT_RAM_06 => X"2F0022A7B5265855E551F77412E7B1EA469064EE2B74E282A8AD6A016B18DAF0",
            INIT_RAM_07 => X"238E2226262CDBA222AA22AA082A60999767C33CC8F6737FBB0E34979081A642",
            INIT_RAM_08 => X"50000081545545544CC2D8AAE26BA5839AC328C2839A0224CCCA22222E022E02",
            INIT_RAM_09 => X"720CB32CB27ECFA178AF48BFFF08AED4A2BA989BC60001555540000455401555",
            INIT_RAM_0A => X"BCCF840EEEEE2CFC2EEF3F213A2A0AEE2288A228A22B8A6E28B87BB4EE2489E2",
            INIT_RAM_0B => X"3FFC6FB923BC30E22B8F9F2BBB046FFFC618867FFBA2A2A2D78E71E71ECC40EC",
            INIT_RAM_0C => X"3FE99E2C0CE8CE8B88FF8F413E280CC0EEEBE6622FEE3FE383BB8A2EFE33EEEF",
            INIT_RAM_0D => X"E2D3FDFC3B84EFA3BDCEFF08FB5328DCBFBF85199F3EE302B4FA0F912E1E334E",
            INIT_RAM_0E => X"E4E2B8BFFEBBEBBC3AE35C0E33E4FB9E00F09C8F933F43BB899B97BB4EED78F9",
            INIT_RAM_0F => X"73F33EE333EE4CF9236374D7CE74FE23FFEFF860CF9E2D3CBEEE333D0CF8CF93",
            INIT_RAM_10 => X"EDD7C8E7433E70E7AE0E33E2333D0388CEF3E33E50FB9FE2B8BFEEFAEFAC3B43",
            INIT_RAM_11 => X"26FFE69A69AAAAA82824A733FC9F33E7F10FC89F7F10FC8B9D3BBB8B5ECEF0CF",
            INIT_RAM_12 => X"DFCAF08CCACEF9A69A69EFE8EE8EF3FA03938BCCF3ABE23F3FABBC432F1310CB",
            INIT_RAM_13 => X"9E203BBE6B02AAB072EAEA2F2880D7C2BFE80E4E22CBCCF3ABE322FCC9A69A6B",
            INIT_RAM_14 => X"2E0808F8C0B88C0B09E28AEC3BCB8ADEE23F3EF1EC0EEE7AEEB0E2B72E2F30F0",
            INIT_RAM_15 => X"8CDD40843C08FEEE25FC84FC9F780A20CC8F927F3C92CBBBBAA7FCB2E6289667",
            INIT_RAM_16 => X"73FBDEDBB6888CD721C80AF2CCCA726EC622FA2F28AEE0B8A232CCB328CCCC8C",
            INIT_RAM_17 => X"204309E24FFFF3CFF3CFF3C3F3CAAAAC4010400440515451545154505450AA03",
            INIT_RAM_18 => X"FFFCE4A21BCC08A33E72CC8ECC3233E8A18C27893AAA8A2AAAAAAA8AAAAAAA3B",
            INIT_RAM_19 => X"43A53E501585400000000000002000000003CF32C30CC3C3008000800002C080",
            INIT_RAM_1A => X"E383E0A48FCF2A2E3B8EE3B808E1B8D5E38E1C832C4CF46999D24084801394FA",
            INIT_RAM_1B => X"21B20CB8529D139021738E38D1F29CB32F298702297B830CB2C8B22FBC8332FF",
            INIT_RAM_1C => X"C0638FBC3F3CA70FCF2A2FBC1B8E3923A0CE0C32CB8C8B22CE38AD79E2FCAE30",
            INIT_RAM_1D => X"170B8EAEAC38C082BFCD3C6CCBD33A233F1BF693F3C9C83272CC9C83272CC91A",
            INIT_RAM_1E => X"CCB123AF3E9B0E74AED1BF3C26E3FECEF2FC070B1C322FEEB2FC0708E88230FC",
            INIT_RAM_1F => X"B7F3C22CBDC32E30FBEAE31D330FC08EEB1F022CFAB233BAA2E1ABCCABFCE3C6",
            INIT_RAM_20 => X"8E9E8FCFCECD38BB45E9EA2FCF32F3F3F3C60BC204BFC23708DAB82B3092D664",
            INIT_RAM_21 => X"2CEB89C38D222551595495955552155113FF5500051451450505155007B0CE9C",
            INIT_RAM_22 => X"F1B4C4B1EEE33C7BBB8E9B54CC4E5FE3A4C3F10E82252554D55549554D554E48",
            INIT_RAM_23 => X"F308CCCFCCCFCC08B17D4B14CE94ACB2E2B2C508EB9D6A59030007FF8EE0BDF2",
            INIT_RAM_24 => X"2B09FFE7424A3A3C4EB0C4F0C722F35F02B080955505528E8CEB0C4F0E48AAF3",
            INIT_RAM_25 => X"61A8EEE74C7C80088C8CB894E332E32E378BC451F34699CDE9B043C31C8B83E0",
            INIT_RAM_26 => X"09CDC6A1A9286ABF48EBD3C313A68ABC2BF0ACA89A1A86A19F1C3AA890618618",
            INIT_RAM_27 => X"CA23AC542B8CAC2A8BEB2922001540008050500505018115054141620505B16F",
            INIT_RAM_28 => X"4C3CC4C2BC6CEB42FEF120BF42E2E27FFC128822E38082E382E2E2FFCE8B5FBF",
            INIT_RAM_29 => X"13F2A3B9AEAE3AB065AAC3CAC2BCA6E2BC3AEF3C4EA8A81EE3A2371E3CC7CEEB",
            INIT_RAM_2A => X"3C67CCCCFBC3FFB3FB8AE3297CFCF329F39CDE316D3CD8B3BA3063B23AB96AC3",
            INIT_RAM_2B => X"AA66F3C4E81E2E2AAB163A67EFF288EB023AC0829AA072C39223F23F25EEE2EF",
            INIT_RAM_2C => X"B0AA234090820B4BA2A53CE332B0A08F3FC42D0FCF28BCD6BCAE0B8AC2B8F313",
            INIT_RAM_2D => X"2093BC0DE96AA9AAA5A3F2FCF2CA82FCF2AAA27A3A3A2CECECBDC1B293150AE1",
            INIT_RAM_2E => X"089CDB9CC3063F2BCFF28B06D780A23EF4C387BBB447C05C060BC48208208208",
            INIT_RAM_2F => X"E3921221280B3BE7BBBC2F0CF9313CFD4B8F04373367EDA131B542237F30BE08",
            INIT_RAM_30 => X"832E4BF1C0B8C1B8FC702CB32DC29307CBF040302C5BF0F3023C1B6F0B828B02",
            INIT_RAM_31 => X"C303F022A3FC5C11C153833C3433FBFB7777767F3D123101E155B8AAC494AAAC",
            INIT_RAM_32 => X"2C0C932A5C8AC8AC83240707C9B1D3F3C8C32C8B2EF0B230CB8363305AE3130F",
            INIT_RAM_33 => X"CCCAF8CB43FE28B5FFC0BCEFBBC8A8C1E74AA52B300CB202CAB323FC322CC023",
            INIT_RAM_34 => X"E7932F8633B38B8BBB42C31BF3CBB48FFCBF8EE0B8288CE3BB8230CAE2F0B4EF",
            INIT_RAM_35 => X"FFFC3FEEE7BBDEEFEEFBBFE38BCB8BBB5E4A928CCBFBFF38B0330D0B88CC3033",
            INIT_RAM_36 => X"D2F3FC4180CC0EEF78300FC222CB8B8AE108C32C164AC9C88FCFF8A7FF2C685C",
            INIT_RAM_37 => X"0ABC6C2BCAAAF763CC3C6C2B4FAF3433428C8C8E88EB8F482F6F1AEAEE70FFEE",
            INIT_RAM_38 => X"FE2E08DFB823332723108ADA0C6AAAAAB1FF38BE2E2AB4FA3C3C2F30B0FCEB02",
            INIT_RAM_39 => X"5D30D38CA13D39E6CEDBABA1202C781EA7BBA828F344F326F320C92548332002",
            INIT_RAM_3A => X"CED3FB7B8AB2AA88BF0820A2FEDCCFFDCDCEDDDC720B822E2EE3883F7F38F228",
            INIT_RAM_3B => X"6AAB5C9B2AF5B2232888BB22C8B2F2CB22CB2CB22CB2C9BDFF4A228B03ABFFFC",
            INIT_RAM_3C => X"CC78CB8870E307D3884F04CB266641528A28A24A28A28929A8AA528928CE9AAA",
            INIT_RAM_3D => X"C28CDF82EC8A231FB9C0B8EE233F4B8599C8A4DCFBE202312FBEC3820F4838E3",
            INIT_RAM_3E => X"E7208CB2AF4A0CBF2C01C4C029997303C0B92B2F3E4A2BFEC2BCA33C48B2BB2E",
            INIT_RAM_3F => X"DFD55C71C7904107DF7DE41041041041F71C71C7DF7DC71E71C7DE71C71D79D4"
        )
        port map (
            DO => sdpb_inst_3_DO_o,
            CLKA => clka,
            CEA => cea,
            RESETA => reseta,
            CLKB => clkb,
            CEB => ceb,
            RESETB => resetb,
            OCE => oce,
            BLKSELA => sdpb_inst_3_BLKSELA_i,
            BLKSELB => sdpb_inst_3_BLKSELB_i,
            ADA => sdpb_inst_3_ADA_i,
            DI => sdpb_inst_3_DI_i,
            ADB => sdpb_inst_3_ADB_i
        );

end Behavioral; --Gowin_SDPB_kernal_8k
