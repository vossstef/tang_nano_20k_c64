--
--Written by GowinSynthesis
--Tool Version "V1.9.9.01"
--Sun May 12 00:47:38 2024

--Source file index table:
--file0 "\/home/vossstef/Dokumente/tang_nano_20k_c64/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\/home/vossstef/Dokumente/tang_nano_20k_c64/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\/home/vossstef/Gowin_V1.9.9.01_linux/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\/home/vossstef/Gowin_V1.9.9.01_linux/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
fKtc7d56dFamvtFDO4O6QlQ/mQChC2vDqB9vvZFQsu07QmbTZwBCbHcSg9c2Qbw2vTp5auoD3b91
VnBrmFIJE7ZO6ixMmp+q2YNrsiA/RSfsNSDEhH0vKQw0LDGQ+LaQpbsQsP38Ywhr5HGWnS7MoDNv
HSwKX9g8mJT7/Q4Lo8iNRCs/QKyWcXytIdWEIsB2yFttuY125pkIy0eVJklfc4fd11sZIxdmgucz
9DaDS1XFvY0Kz34P5/p6mjfi3PbE+sys5c+FAVy7ctopbtMai24WShkPhMkbUDM6WWXWU74ohBRx
wu/SC8lLKIqFNhuwDpfDWYbmTo6930i3iSJX9w==

`protect encoding=(enctype="base64", line_length=76, bytes=15648)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
J7OqTEMA9RykudhBJQCJM+4vS4/K1RGZOF0Pk7lbMS3FUL2d3QM1NCi+Z0Sal8kuPU8Dxug1AABP
BWicpg9wMh5NT1silzRp53+V/ENqIXDHSFURZR08gdBocwfCNe3idKO0aEcbd7N4r6ZA2OJ9HnQJ
YzNjA4UZnR4S1oj/OxEDwgHlN7Rx+bA2MPhCK4Z7JWmkeRlYUs4IxGYBegoxc28AHLfcQiFb58f2
762lA1e66mFp1H0nEAjIFhfd8EsK1XGaK5zlgj7K1aN0kmGi3p8zijIsUsj0y1qTuzkKJ1suAbJf
JofCGdWFq1RzcLQdr13ZaiQhAY39ikv+CMoetKUzLyL3HozsiqU+TtJ+HAxEp5uq5bQnREj8I3uk
Wq6hYWxr0xZpFG+ZftzArPkGzrIYzyxpx7phNWSt10dYfPeeggThSGAigRAV97QgqkhAn8V8PXks
deKqRpF59sgMc9YxKPUd4g9rnF0mn+8uCo4cWdu8lSK7ZXsMDOVblvkScyR+xbqKNQkHIrgvSH8A
g65lB/5/xoSPWHi9C05eeMQ+uV7E7kl7mBsifZsiHnY6E8LisOX0yXmJoHZW5bzfdZRNYqrOF0qG
3PiEQx5YFJB7mHmi4dkuPe12YQhNyQNMsV+doW8v2lsKef3llqzt/vnVbZcuK/Z3STSc+70zRQ15
7HCXdFZnEQCQYe0qpi/n4ufI6cdpMbTWJL3Ryocr017b0fgp4a3FzJA22G64MGnwkUBvznF64red
NGkIrLgRozpUrTamfHjAeOsMnzyxVyE8oUmWH6SP+9eV3OQAk2+RWQUGkKbLdbO4N9k6e7SfIBJH
j3UOlV7SJvhODAxHJqp3twDjzdxSr0QNqbfJFy81wdlVinbrIigLrbE+nqnQQLlWNdpnZcdIzJZP
gJnBjpEjj8IznGpgeCV8kjfqPGsH5yAvlVXgjGTGlnjwaRu25Y5yoIFlHanNymS8Wbe++Gna6GWP
8B86ZUS92bNn0b1OVXju/EmayQMM+qliBy4BFa6+8PkcVsRzEXiUMI1m7SZhlEJ+BLeZszlztpwa
tz5MCWI86ld74zEkKVGZdiPnjvQgj9gfwH3Olq1Ug0TcLKIyzmGvYY1FdE1C/wzoqkf2cZzEw7z0
+SqvwE97/EdJBNVoLeului+zBk3trfsgGK1eIFnjLvKuXObhJD3sibLjzs1CUW1sRP8tuaK2yHbl
aLM9BOBU7XRqP8K1MfCt5GhwrMc6c8/4B+/yMBIYd2dHDR1fayCqS95NVZSmcjfI8EKptwYazAQf
lJulXOP7NZ6aUr1Hvx/ygNuGCiLKRg1Tk6ozg0JZBR+aLJzpfHS5UoNWFInJAxzmxfukKsqF3gA4
DayO9aKnF/YjuYearnO4JjIYH5MGSMMAjcZFo+uW4ujno0ylNqpuoazvrT5etC7G4RsOC2sJSQ6W
Vv5aZcZmklRQvB+B9tjpaedftfxizpLE+XJKUccTxJI9OqfYFwsUoagBskp9Yu4NbRB9V1qjYmPS
/mcj3pDh+xc4e6Qrn+bRJtzkWQMRkKmtD8mN87XPY17Up2FXBmad/JUr5kQxQLApUQDY3BdvRBN1
LKEbmVelVIMwU6OISf84/2P9nrLdqH6zLyIzr1eAhDrRlt4Eggly7RAQ0zzRdc/pPiI/OoHbB9n7
3kh69YnO5FuuUpwkflpe4IGpTEHCIXs/AaCoeeTUIxvsWMKo52f0MbH/Uq1vaOCv8B76LnAwVN1n
xTYATBdZ2E8KpFt2u/oH2Mu2+fowsV8tIK/tEyoIS5SKgrnkF8UxbKEhClYlYCU+jDFgu9gzoOO+
S1C8d8fMHRX5pJM3MpudDe2Cc6E1G1vPqm28phgDsZArbnz3iSBfkn60EzqQiVb0JW4ayCOvDvSX
cvDCa+GCieO+7zbYavrQ9hc1f+dtG0L5WLUiC2yDLaHcL12Abgvwb2CxgIgQKdUFhH+Vr7uoJ7NC
md2DNFCbd1zc2dpK5IpYRrl9P3xGIkKVacVeBmFhRl0dqroZtbbLGF/iEvZbULqNNmTpyl53z7XS
KEUTs+pe36DxwEV6TzIq8+m0qMlXCLJsllBcQ16XUzPlTjLEGasRkSZqVfiefoHB+hj2jzsoEU9p
OI//j+Cirgb3jwL/hkZaEIndAS4FkkBcpHvNbvLkg/R8LdV0nkOgQHGeG+o1hG95aoxHanD6BEOU
yOuYboqObCT9eJRhzTC+OsKEy7fYCRKIHxAU7RJZgQpGzStbgF714tJLhlGMHFeeiC55q0paPDY/
vZnn4WYe2vgapcgP0riPgZfU1FZF7WO2s05+ZIdzrROITIqSTLglDbuVe3ilXXyRcEVZrgPLcIY/
usuzX4F8VMY8d9FaJ18o7/DS1C3m3RXwWti9pUWlo/ZwmxDRpX6Dg/MpsqRGO+OabzqK81fe6GWe
fxDm5qe9ceEzkblri0v3jwUYGIdmRwBCanIYOGB+P0PTOGJrA3Gu/mQ5Lhb0fsE/Bxa9SJm4Dkss
WOMmAz3wPJdKPUUo9W7nssWrphbqZb51h4VBq0M5ILlwrKdJ5FEeWJlihiVd0dyBWVDgfOF+KJJr
BoFbtwZBpZ+oP9MGWlNN8GKp8EUOyKWlLL2FczyBuOflo+uv1ygT7E40lk1nt7iVVmugCEooH48s
K2Vn0jVONA5VNAaeqc4xaakcr64q/lz4kb1NWcE45jgzC/vV41lgjevDP6V9CE49hWCzwGdufSno
Q9bD1EOK1umYM0uueI/VbpnND9ZY2o9lCWebeEeLn5GxA0IIlYqvUhULvRDPdqX/HfIbp2f+xDOn
plg+VA5nUIkr8kDyNwiVPMU5F6jMzzw+g1R50BpsKDsX6jmz/FJU8mytSbgPElCrv0t6U/S8uvPE
zB1QVIshzD4hf5gjlOc6TkqnSnePgViFZwiX6PGJOM9oT5mMZsWMk/NS6mcg7pPlV0sa6zbyQPNO
PmYnKrkx1wQH7pxkvtqDI7KFrOLxi/Xh1WQ0pc/C8WFk0pOKeHGN8xabOH/xBPsy9/VmlGDVfNEE
X0kVQkLpjYQLqWWC6j7AxHvq0tbkd5GmCeAdX9awAlmYPDiVzjFrvVD4NFQDZmqGRviB2GrFxd5z
vBBlvMFsRpLC2QbbrEeTzgZaSrmK5V754aCJQuB4ceGTclcxU3vCAqZVHskj+W3JHWVrpWWmbQEx
JthHZFWOCNUJS+AOMB6Hd+XksxcxjNwugOcm+DhQNDmvvBKIQdL+wOFcbi9aVM+DahAZX7x/xE9q
Ev3PMln6vfJS6YMz/QRhKFXEaxPdAlAncMbIFPVcBSVaCyZqkpUBykQU9SZ2rJ02sR/zVkMyUrqe
U8WrGGllQiFAdZ0FqlDb8Hy3mvVSrN3Zt98NVnijlG+Q/Ycy4oNADmprsXU9HoCxmiKEPe96QvaW
60tJJFTCPvn16ubIDNkdbOAhRJE67PREwCOycWFg8gAa5rVpkUqDJTzLgTDsrQFjq6S2HO4YOSCT
eTzjDbmpVH9AftQMywD4EWoB2b+voXH94Ww69xBs1S3uz94H207qvd4yJpH6D/Da0oHTAZt8aaQ7
V+PWDcTw9aQXUlkKbA8YlXHlEdX95FE7hP4Scld5S4vRZKcYyEXuqA2uHAc1GVvv3HhthGxW9lAG
gGk/SIYOmJMvMXStmT3+GdeayM+K9LsB/DiIiJuEaSwgXodL8vDgCsW+eXbsk0CfgIEQefykDzBZ
MHyFoTch6v8T755h+YKwqBO9EdZtY/vpKZXZm8tV0sBGZFtiVaockEVP8T5oOrij3FNlk1wp/clU
w/2bjTK3gHNcpwhn6zvjbX6TxX3dFGBVZdtSMHZtf7xFIlONdNjJPzyWkVmQtYqetA33jTfQzxqF
nXSgzN+L/xBRrNVu+h/Jq7cVEUvFvlWkHAOhXi8Gw3aU8OmG0ZVlJSGkCIl4rHmNjgkJr7q/PQjQ
PqHg67CfXCF5nlgX1FF4MeIGmedlmG9eX9nUGXPd53csB3i7Gfe8asrem9iCQfcyw8FudP8lkTvm
eOMec4+o7XC40NjFxZv1IDNMlDR2Rv7OzDPyxkoLM+uSr/32qLhbT+s0M5DB4X86xFoV6TJ9Q5Rp
jHpIhMLmCfcDiClXBQKAyel5fn29eoP/xRGEqVvqhkoZ9tkgFq0SqHKD8cEROjMFtYn8oDJYgeJt
ffOKQCaKGBPxfXaLq2vH2+N3xzEDfKOqSmKS9YJfojv0bPTJTHuyvcA28M+iHyhJEg1f3iPgo8wG
R5UR4vmrIkvrO/lj61TmBgHl6COt24Gu09FfQFUrmAU9lcZQ0gUyBeaqahXpNBDPQzVA944/w9kJ
qyuNIw7O1B5pA82sff4nmlnyTUMI2dMjX5b/HnQXGK8EuUDwQEUW1re59ElKgvIoAKvoIIy+sEV/
W+srKIe87XtMmXLCIaC1kgs4agsT8XMR/oTF1y4modygfLA3b+pREAsslwZ30ACi4assydCDAoAD
OPxkuencAnOUc1LSeoQApwsiJ7Z9g8BfA4O/jpN3gfS+5MkT0gWbmuPlLyjJ5wyzOF4XWcFSqRX5
5cPKcNTDhPPcFQK/3hM8NlpijdUwIvpSKYBuhTQsZpmFKBAPz3o7ABfxV4zGVQRbeOfRp6LGbf4J
52EhhlTt33Ja9PcfonNH8PuNfruu9HUMcoflwEAquh7BmczwL861T/rNv96H59LayVVFMWj16blb
M5zYTH5OfVqOYmYLDkqHxzDqeMswlpxZTVPlwexJfyc6MPV6IDTMAb5NHBdAqzLO3S5h8wXq3BkZ
6u1FxGK/qckvrAwD2goMjxmlQ6vyhli9lvqxpAtzliPlfbeqYRDdkweURi6Q85l3Zcp4EEDtaC/S
2trGKrd/zZcStvacBU8Z6jWaED7td5+p0Uoy8BpdGbnB0zcTaZngaZmojcIpzl/Fpcw+4RTKbz4q
0hkACA398jrk9aB6KH5317++pHypt6DHXk2HxdxZYvEdk421FUXYe3+PyaqZzg7xjOnAmRzCvbh0
sZ+rnvu8ICNMnwOF4XY2h6FN0NH3qvcxYwKsBCUWLF2Qtl5KDVbffZ1vrQN3bko8ruFpruWOSDIT
z+yMFcywAsZ9b0/5AATe86aoSqzAPU/Mczc2/hioiCoCHXhziS+H5TxOqTyIp/ZCkkqU/KWinI5R
TV6Ir8/c52/4hB4jAlzEpqqinrI5TU07/1YEkFxcaIKlqiJJ2pGw/7Ckkoz5PeC1DuC59RWniPp/
bzK/BrU+sRxY4gQ6tDONOSwiCLQsbBNM0Jq+7hwGgwd0AmJnZpD6gBHcd2uGdZ5Aajth+1+7Kz2L
DkKUf150D++XVeWSjOYf9PFnqFtGAGfLz7FISXnkmcYd78+dHjH5TZjZyLednO3MUI7JFDYY5J3C
XMsfsZt90pSuZyFO4Si7ZXZGhG9x1gKO74e3ptRnzb/Zl9ANisjxNSStwDJJxD9lqwYMulfg9xQV
RJeLWoyb/vPmaEbiHeY5ZFNMoo7wCte0AoZKgc1BmzuXBiSb+F787KsVvEvb2//cHHYuPkG2S31V
DVznK6gSuiZabmG8I6w2Mp6BgFfgoT5nZofAexDjjaHUvwAdTrI7Ng/FDdg+B3q8XptYNVUG48pD
GqgGiTv8R63zuDNuxAlLu7/BatJchissyPNWHK+n/8rXg3hoUz1rM/u7nyctjEo+jpU3wy8MUakm
rItuDRS4aGHNrW67pQAbng5Se+vP73/ofDBSSxIV1/GbUUtT9hjnPKgi3zV7tQNZZrdpIXfcmcwS
35go6s3Gd/2WVW+/X9bgPqHdbcR3X7UVSSnm7/n+Qz1o9xu9suZxy6wBuF4K9y58dGP93nKZ01T5
P1yRhS3wiovs6cJZOzj3MsEB4dsrPWFQ8fOeZ2vT9nlCPSxX6H7tXS+NRJrfRtO323wiIoo7uM7/
SlV3eF5JcBz7kEi7w1gfZgvYaoOXBmUQWaimv71hvILdCy6mV0IbYnjsUF8pm47rplr1YZaUHu4p
HztUg4V/tq4uItGYkzZb809d5z07928Lcp2QRxbBHiDMi+EIRN0xtRrKs+1tHolUQtS21UCcimVa
D3I/wtkCcHpuyF/bejlmMkMzCbDZdG3diHlinZFaVK9TPiw8gNVbWRthXofDtKqpI0bLR2uMTzQ4
iQd+Mb0ShoiBwgfYtZHUL7Iva8hwItPsM9NUDGmvdmowpH2GzR0Y2A0wcMxIzXL7PYVIaZhVOw4f
Kf0dwqiiS7LFbkn+cBT9+v0bGDgBeQgnFOqhMqW8wB9wZ5uvGGBMAML3JAuV6TK8oIkOLe5xXv8p
Ffnl2e3smHt8ovPBt/UWFFp0+MwGwnfSIgp53oGtQGZn/aL6VDVtlcyZQRpCgiRjQdj48iXImRt+
lrKy2YNi3+lyBu/kKZ6K7SQPx8mQhddR0Az8/l9tQAXLE+pJ28oD0PDTm2WTTeIn91wblYcCST13
+bx4vXkL91XJjLLtsQSeiT625NRsGBgxC58yoXXWRDRKeI6ymrZ8riEZY+DzQvkKSUyj3YkDqIuF
usmVDW1qhpjZN/emsvRfGlUJxn+Kd2qDowjnXbZxx+IB3tSAWJLIuM2aHKEMYnMx8R3UM3gOvGtc
hfVndel0a4WMv+uiukKOYroHBPuNgU4nzePyUdiScXz50zGU/Mrsa3wXpXDiVueFHwnElrL2qxRy
rlWPaKzL0okhhr9rBVfBUdbY60JgFL8ZGCPyptA0nTUW1UYWeaSq42PB/m0osz5FxtzqlbeBpUH8
jlemv32eYqjGFDheybndNyyKr/DZbHyQsxUtPa4+ktGO/dw1WxJXk5d9mbgIhlJb78tEjXL5c06B
S7zod3J/iMbYR9k+BiHRaZAl3bU1u2df+96eeEZsX+5yD2SqvMYlCor33Cjy5eE6itPTd81/BgoX
GrA06WLtCBNLbLAe/XjNd9ahX6fpdjVaK6e4qT+wOvXQ5HkpAhMdKb+H+ppaTlK5unHLD3fbMfvQ
uxi8OKwf6Y9sxBlo70eQm604G6dphM06g1ocj2KnZSWYnbY+6A/akWf+RtjQcInMaaZgyvL38Yb7
wVYFGYQ0mFHcDOGwM3UGjs7lzzoSU3/iU/ReCTDqCOhr+P8m5O0m76yFBoN7QNjEJhhaT1PkzkVH
HZ9G8Lv1qnt3YloDkW925WJqSg4GT4NP76j0RknTtxttYOj7+VZNP5VbB1JAPaVfqChU78pfhg0G
gDCduncWm9xOMp7jOSHl8AkbD5yig87Nsmjt2k7z0Z8W3jiVDrF+KOJujXAM/bM3Mi4OcX7R2WzR
1u/NUr7DA47QCeVQZdc7yyT2D4XhBDblmrIiMA4ITVPJNF5lv9F5QIjjAH6FFuvSF+KYx/zFWvdD
+5xf/5DGSlikxPQlbd8M3yQE3mNytAsxJDxXsuoCnJ3BnRmHL5ufHuYoJMtL3V5/KDQkRFBKLsfz
SSoCbughLjIHq8VtvU8Cuv8J1YuA4DaMZ/0fAyDLEA6tVo0oNDmOgYeuMeOsoIsdFvxzSKTpWh+Z
yZn0BrGshJM/ZYEB+czeXLAdWTuoMDNOanTT86SHdOUuJIrUXaqjW1U+4d4Ovv7XYBPr2P0xL3hV
+WzfFlVoQ0XYsmH3Z0jAzUcp8flPGO5bO4ScA4/IRZEOjwulNqfOHR+3m9zlRefDNyAtjQJDEy7K
tVdv95k+6p4ozHYeizBlog3VZz2eSxIWN4SrAZBRkHJwHHp0ZFIsdV4CpLXuyAPjV+UYdNZdBlMH
ETCMYaBzZVsP468Ao8pWJmX57Hs/tdPaxEOJ8Y/ub5NwXMk7GLzxr0WOvmzoXZmd0kVEIeUFfHiF
oc0buUt9joMDFdU+uMm2FC4sou1qkVk6YD3isBQwYI/pnjclE7qhOnYLZCQZI7iyIJGNjbvMWnfG
QEyc3t/vvIAsW3EZCYSF/nEptYlXmDa/1siL3bX0402ZIL6YUNNc6RTTpA2R52A3zQaCqh+8QTW3
t4lkJdfCOcamS1C6xfPPtbig54KHabcwj/1TVy36/ifF+cosq51p4xFVStxGvKVRmPg9rYu4Y/ob
W3fzYqIf5JwLERqyjb0gFWSW+Xups2gFvjQvYoJ6tIU2Dw/TRYDgcamQDRkCLoC7J9h6MJG6rDx+
HApc6NvzDqK6QnFU9AkJ9AVe4hGmtZdl6JFGXQLovu0QPiQFqXfYCnJvjUh7BOJipqCg8cLimT43
guDACxVaSiHGoFMMIRYeWVqM/XmZpTJ2D0CSA4dUYUV/KWBN9WpD6XvdYMYHSBPYZLkxiPaadS8z
gxcqhhJxTVVzILxVooU0iaMeTukWoIjJIMmZhjXvntqFxxXo0xQ/aLsInrOXLIXwuYHBc0ffTlIW
MhCxVo/sSZO4WK6L2mFWlJcpLJ5N/TyQvXHoGL1z8Q09v9Q1BWHdGjQhUtK9MFCVmDLYL/PunsvY
roThYZWZtMGaeA2js4ijyXm4o8DD8FdQ/bcrzIWzcBfIGEeUBAUQff1fBCOkH+iV2YJAMpxBPiLh
A48Tg2wb7DLSsQsZtj3SioRlYivpMZOY/Ud4nnLgemRz7oSQiI+qb7/uvVoxrHKTUQQ29qqh8YW4
8DIwQvMvmYOEPmJ+SdEC2ea0xt4VqEvv5kixfswJ9K2lhQanfIVTTunmA3BRbAeLOCwk+4ntX8yY
szSb02RVsZevZd/pv4urYyooMP2z/y41HKSeW0/D2gfxfy2e3vqzLUXzOd1rHsP7Pr2GOpGwaAsx
eNIBhrnYNwgjj5MVkzw2dH0iIsqBx3GtLseobvhzODXibYTqWWc2BvZh1DCh0fMH8+w181MsMG15
8DABjBKVPQHrltRidXM+bj2rEqP2wN7gFrIgaQBR9fEeswh7T2dlnFuWl3ZINMGGtL7jpQDAWLON
eFz1Bp3rXN9wEU1Bx+l8Vt2om+TXQZ37oP9owvGcSqj+xhEYAHaUOGf5WVrzy2ZNWt65U2NvtDxw
k67EB/voAmvxib8ewQH+YIHNiXq5Z0OWJhotby4hM013PC/gD5taaYbUn/cQ5GXhGFW5aVQRis24
W6EUn6SL+mNwRivcq2RpNTpXmUxNuKUUThMWmS2Fqx6urSRdXkTgaiuZbf1usbfHngIxusQ2dd4K
jYnT17gw0LPLCPBXDuskKywWyoaWlJHYBk5sgdwjrpEOkqhaiv5U2k4M5ufvdjvee7IbzwQZkPKK
ORyk4xjkf1v8qhFRYoRDAaau3Ht/VN+e/46A88u0D6jvY8lESpDXN95crXRLKDTYeXn+N1pllcCs
qoeWxBkepnObwN1zByDXFKJcZbmshTrMsh6/E8g5SaM4z5Uq38JTciPlHFGyIIQPXIgwRsEBUChf
qVLLaH4JqnWXPgzr9pvMOYbGN2yGIDvuT82CvjIc/Mgjo7sSynM9S4qo46Xf03lK3dmZ4WrewvYc
mo5fQOHSe/+TemXaBWFKfxXObMf7j0OYTOW19JqjD1/6lY8VaLU2jK35R7uDD5NeFXXMpJRHsiLS
AhFv0MEDb1jDDSQPW8HCUhMsnGiDAdrsUagRbEHrQCWbbs9essSQqM6ltdn6tuih7ufDWIV9k/Nk
66vgglGer/zbjG5B4CFLzb+z4bDBSDZhMt4LGZlX3x0Api62Me1g4KAA5u5wONcaPaLqBHS1oGBA
cWeq0lhIUE0UMcZRc8+Xsq+h+0XmcfBkd6JYGO+IIOEWiNJc6JXh9EvQbLI8+xokEfKVKtq7IIrr
ZAmn+s3I6ohgVhW8WBKzB3n3A5ndpfoxfDvTSI5e3y/hpxCUNbtxwN83BhsaBIgTdn4sI2WVm/QZ
ZUgAS+tIC47uXZbbEM0ILADuR453rCwd3prM61gIDl6wa5tXD0WlsKr3w5/7Y7ltcjJQih03LkqT
Dl/pLfX8BVIKb+9/dG52Bw5FzbtGU18afIFG5hlJa78vIYzOKr2dVwAy5BQ628JZ3ix3oyQANmFm
xiAHpcGDIXsrriDg7B0ZzLSBxZC6rRI50+BhPdLLN0X1C2xQf2Ww0k5ITalEtHF4o3H3axtlRfth
cvvBYhnvKAkP3/5cDe4aMPUKIP7buX1fI86okxCec7lIBBG8tV+bm+IdeZRVRzw90sTD2X0mUTye
/5UkJqRrEaJFzoSSWlrcv1wyFpEPPqfSdsKPbZohMPKTzxtk4zXw48C9gPpzQI3Cdz3hyfpSf/Ok
mJvIusL59x76t+duG/tQQ9WiBrc7PhRyrDy3A7DZMCDb7cqdrZYWSz4U/xQio9dGhV69lXMI7RJN
L+rTL3o2/JMCUJwWtQH/y7W+QrEL9I6ocLSZUlQRAcBq0yOeDv3JC2kUC7g6yLq7HlRGUxGAvTNf
sZZpppkU3b1TDdvG5nAaSIK8RQmkwydEo7BbQcwgREmrHKh+FvsVnCfqWiWutfWM70cwE5TWFp2k
7TDt4LO0MTG4Vm6MsF0HzffA5hkSiRsEIS4jTuClibbZyS7d8AWCsYGCEV5uK3mrI9CXQoj26hP8
6UTJpAPJ4L/ieZVEi7DLpjeMIgp1rA6M9MkDSyxscWnqhu7dRjyNDrSKbPW2UZAe1/fQRL8hfYhG
jxXlO+bOyBxkKfN9PxQ0ZDXYpbpEGZWVkrrZ1wwjTEtsbLl4vSoZOguT5F0yZMIn8YGKtrBtuLbs
BoOzW5vB3D2X3fXgzYmphkBprX3hVQfZAsQ0T21qmFsSBvemYcyWwfYH7EdckOBARGAo42V1snWt
zep4BOxxi8AeJbP2P11OsFNMXRTwqdP7hWpk3/WS0IkZb6qOMp58F6KQ8S2UQR53WJlpwcpKsAb2
xG7NB3KrBqWEJkOP6XXYh2Wo+Mr4nmLSuC6yptLT4vUPB3aVg5CfzMhRZjWUMjuJi43NDch8RuJK
ZlmXoxQMCLSvFnH9Mn3oOFAbGD3D+N03T3jGnsMsjW1B09vberybUeQpm4dkXhi2lxE8dgsueoHw
Y+jd33s70tEuIQUSgPkGw8QLgfl6ouajrN7SYjk7P2zGnRaMCHf2N1GO5f7PuCJ/vf0Gr5qt7ruK
2NDtmDTeW8RkaC8sHyMHCu2Vh/UIAI4rXE+Aw0dExz4qbRq+UA59njMJSdQTI4kD696gwSqFe76E
ueZv0BfkLybzfnhRHZJlIqRD7Wy/2757+r7up18es0wwCji7+ECxxHBBLYVBPoDCVaHLi7GEdfuJ
IVEWQh/xOJ3llh8q8stkMNpkyDUfpTzMppx3Kz9bm4Pv1onTelqzoVpOY76atvy0dMNMOCXJ0+Qm
2tWbiI4ZL33clPxjBs+Q/IZiJrA2JTzaOhv2eudzVOL8diX5bFcMTUXXDnM1ubsxC5lffn5wI3sk
rzbH6nmSgYSL348AgBYiINHoZZ0OkWKWrUpCqxaF2x+6512dgYFAupEjUxScqV0H+A1sR6VHbgVG
XTH5/7GmgBgIFMTV8djt8Nw6nZmBuhp47UtEm8xX+/P20AupBEAxrK71EBag/3rIDK+YYRa2WW3Q
DUSQVxdAC4qP31HyB3+68Cyz9KGg3zIjl8wM93UT7zpEknHdTdDJstY6N5KSF2+xal/ZhvHdl4Pf
8FDTml5odNSg50Ry6D2iSsb0QNBAdpcklCsRDyIgk2uikkE344/F3NWbXAXlBJO7yGkh6zeMd37h
BHAkzHzykDSWGB56vE7p1seKVtzs/iGEeifUFp9jpUWNlCL3Hyno06zwjgpeaO8EofrshoHzPoCG
nccefQ/Qkn+l9PMYWkUVniGbzYSdEWhaFmfFJ0rGDDELzpKHogyWjga9xaTvgq0n1IhO3zsMGf4I
wHU8FNG3OvKGMjHJ9ahAGh0EPJY1Bzut9kllWs1orNYok1KlX+eHvVBwzhR+wagKzKamomSkXj7l
CXvtiSvTWLBckA/VOKfgRSqifQ1HRHU3RQKH/6/kYYJCe8B+W36vmyO+EhKJsPjmGk0kRlYO1iQH
xbySq9AEVFb6f348/QTkBlUurv38+fLIJ1LWEk/E99zqoNSoNTjZlH8PHdoC0uVEqkfcKiqSJwss
snGPP2DL2gc3rm3W2l+TPLTK0sH+zvBAfOqpdgHk5nPvEFSNixbnOqd3QhTFJg6BNeyNQMLf3yWr
8IAVD1fD5kQVpvaitWI3y/tuFdyvsbbhIeUCGfumhuE42AtuB0cyweFq2xSdQRmgwiXqcrFR3mpJ
5PQmKov16dOkSYeuMmmEbKye6siJdl9L+zShbti1fmFBcUe+PvS47y+vj0TzmGz+QSsr430MuE7M
Vp4Lcm4CQdvgLbORBBpMgYGiAB79bNhCoxJ4/gist+7aG33M+2FDtkB5JhCi8pCAc+wppbtWYc9Z
+Zvnlo6aEPIHA4bno385QeveIinuZvFjoHD9GOsETsn2dULXfS1ckd1/GNe4W7iOlRWIlkIqTbm9
oV4yH7srgDCrFOlFta8rPBApFQN2ccy0H8fwFE+qlbsvVmCrRBwrYksbLy3/Ofb0PVOxbGyF2RB9
wyYxvz9hxFS6a60T0dKZjKvUrvSu384OID3L5PeR8dImWStez5COQy3EhQmKK7M2/2MGNN9OwNB9
w2cVwtz/LRYxvVNzvoRk7OXKURL9hoj87qmu7PhcFRraJD4I7mBKyjqoSBA6Ikup6goaFNbmtTcM
COp9NQg3LFMhChweMIbaLgg1QByDkzLj4mfahysf8vhZaOxWXYlh0rKoOwvLhds/F3ErjQ5T9DZs
cXpceXr2fXuDYLJFa06MOC/aIHZnCxcG80D+2HEGlkx+VgYew0oZmDvZ22aJkHW1pfvo8xL1goYg
EnMFiY/v24YXz8jWQ7quAHPc6a/n3XDd/ZwsGp8OP7O0ymrL8La2h5PPjYZRO6rE82obruw9/Dou
y/AijjGdj5gdkUVLSIjYypjqw5T4RbHhcMlURH/lu0fQGe8KswBWoFASR+Guf7kUEyy6m7cSQQDR
pdLwaHwsfSzY+e5sw6IgLNNE4WnmEVPE7E/4alSlXUr6n+N+c3WZTTvlW1uzDyeMI7qxoFbGE5nW
04KjEjJ5UyBKbpT9kHngBUehi3Q2ZuYY4R8yypeIB4a5z5sltCxwyp1xoZQYwiE/ToQ3SRRz7pcZ
BUKtDzbxkweG+nGDGhfJ948ww/HhAX39QdcLnfZoUmkUVh1NdcYShHcWpwawZu+Edof8lgVr+G6A
WkHC7k3VlOVTsofARAIPEG10lFUqp8hCq6On3Hc2EG1rwI1Ce+QVESPUqtW5wSIVfEJ8AnJGEN0p
aYbISUgbqn/PVFE4VC0zG5Qlt5SqoBEIzt+CR2Lnzi1h2os9IOioLlQRZmTS+2hPRPsAQJq/avjH
w4DXQV0YOItha7EKw2tNGUL65/IEXmvCx3c6ubK5cW+15m+knPvrwr+ST51iXZ7fbZdp+SgP++Hz
1bcLdW3x+P1PNsBFiPKvI4n4RgXLUEcuYuoFl6VuvMB+7P5ZCfLb8TJaXLFd2nmEjnKndZWpPdFZ
vGddy6Oq+yEp1zzQsw5hd2vC9QxDPLaTivegxvN+uuF+us342OXyI7/hBiWhbNynMBwORzl9bnwu
47abHOgFHdMgX2wtR1QHVfT/vy7X07wj/RUokLyY6sRMoGAHoU4zw30f+uSMB49FecOv2LdnAKg3
KRUSA9BxpdHhL7vqEjPmbMBCn2SEEYYVlqlzdzVkT+svr19TR+Fp2+zs79wvmKtsuam6zxzYqZS+
XoJTKqhTQHKO9X/ljPsgT5oxuJGVAHkaAhBf9X5OJ+Atkx4nA3QgtBfHs0LDoRHp5b1Q69STeow/
Nr+EWAjkNNvRguDtq7frEdXW30ZBacw/DouTfMDcEObk+xJMJzN31LjR/ffXON1vKYKwa5Zz8zTt
pggCITCCmV/7bbPDpVphKXfBDR/cRUdM1POJ8Mf9gNczTZOiKtUapv6Ipy3Q5UfuaMBtWMda5EFb
Kad5st8o1vqs46SGq9It0wuI+1ctD3bwGQUCrvakZ1Vtn3Zxdm8OUIE4hf/nRiktGEjG4y3WCE6m
eK3Xlw2clfah2z4fBInJMpQYOIydCs6AT8HngDVnS5GEJADXsUOO4NcbgQ0fTZsKYPyy5OCOfVAs
nOXgYp903DEFEKYiXB/4iU39hYmfot/e5AJMk3QXqVgkMMoT+hU7scI9/D11Gqm0hyUozlos+NFg
trT/0RGT+DgqbUI6KR0nQ9onSw3ajW7XCP+LrztaEHzr41uOifsQ0Aex65gc5nmvlbWAIpiCyNpq
FPs0ckGMFLaDazZix6n1LnLR9j7rWA9sWpCEkLmpgV8Kk1g6zkrbHmf4pqRDWLCt4csp1+E7el29
sp9zFxwIzA1q9G3JHc2pttQ2w5m5ErOVdxPSxtcOH4j9fyjykZWbUs5I381mNUwyF4vUXUYpGZSN
OeYVNV/+0cvuhht3516h3UnHez8SPTu9MO6oxJjI+CQChEDxfILWItR1moOj/RkshVdO6PaCAebu
6l2tmh4jerBjDLxdDYEOh/xdYLP2GXlBFTSsoTtSH+T/WrL4Ao2/Nqc1SRSZa9WUdD05KpFSJ9ih
aUwELNI7hxsmBW89ObvpPToMrWPtt5Yny7vqgqBz/k+wvf2MPct0O7M7CixdHMJBI1mT3yKG7I6p
UGBcRn2wrj2oiBOfWb9PTS+ABDtfNVCDOZiLxl47/Zf1Rs1uVSnIRJnaYJdyLYQsBo2w/6On+B3K
tfEdr3RdMuiTOctTk7JojUmjvFovgNCvWOR1pUlK11msAc7+jCqExJzdxAHsPKrFbqv4jnAWuh9p
jSJeEoVh6FuwZ+twSeh/EYxScGmh4P/zoLNnnDZjfXq6Uz4M+nSJurHFcKrla2p6Q3xFs/xcnXo2
QVPe7kicAAZbPAXwg6aS8uAmxRMv5UM09KrQISQ/9sx0wIlacs3+GMaxHVf9r59ZLa+a8woGm+rq
9AonTEl3URMUm2Z2xkPGfVnBV3qsZ8D5XvKGFWd9rki6WbaQnJay+YAPEIWNGT3ew5S11HmLwySI
ZcHQWlvIwn3YKReogx1IN/s3mIvjSHM4K5a3L0gpzAAELRkim7cDqZbN8dehzmn7Iflarm+T8xVk
X7E09J8COXuXFIZCt2eVxEEVOecOuCs5NJMDZmAR9Jrb3iOzShChsZxAcLLid5Mv9QKr8gGc9ZqN
0PIRwsVZfkPoMuSiM8v4ucTR/ofGmgoBqGp9P/B2w0+gzuBuowwSdQdpxD2QAhdG3CAJJmTsPYaI
UJ4tgCOXwdHqVnbPl4epeUdMhYkCotFc59gTNP9/VNY5O0uSCk00GwLZcWGJBUMRDICPaJbhwfuH
vmKyACOaSIbQyjKq8uuet5ySJllZq65bSrci0A5ruhR/dY2NCvIN/qy0ZXoe3GEUuRhTpxZOlI9p
3W3xHz8u90ZIrmUmqJ4KSexhCnKg2mWTD/PRVlalSX96uiRkLrFqS5HZfOfBHDAJfT+pSlP0cguS
vYvdHmHowXK0SgKp2bcjLrK9+XtPplSPFEqBHpc8448kP9NWSqJhrx17JQmyowngcTs7MFmgv7Bi
Np7CMrYH8EqJq2vaIOTjTGiwTEG+42tLid28cF9B2aibf6tGaKWmrZZDfxnAJh7aOG2/duqGnYuh
t/0sg302p3m4DTx3K1rCGaytEQh8tDpE95b4qSAb04hNgXGd53E73mNGrWkhSuyc3jgj/SZKGlDz
n84hxbttOpkVpsU5U4YCg6CgmGK2jrJukorgwpvHlVQj2AKaTGQUPYw78dGlHTy2iYP6VGZuwYlF
S/csseATQ34z60r0n9XWyCkPUMCaNU7gvhqVMOeTGnPJmueZ4DxvpX0Ft6JoAmLRjT1yxgrDPdyg
sCzkIa2zDtgdBZyuUjpCawU+Trxao4KPiG7xOCk8/bIgWoB5tPKSOsvJojgkiW7hYYm/mNRRSF8b
JeqLBGCtjinzaNxTGkDRy6jKRid/PDERzro2tHLu+lcTVTO0XF39Sqa/KlrCcgP2OZcmByIvefbR
9C9F4lEixVjD4xNCQMcvexBxxgdG+ZU140X7Qn3YpGLtPdtCubUkkQk3SXcpZAhtOzD+kvUlrIq/
WUp3ZMpol82d57XVXA9/+p/dr6tpJQNFpouhqRThzU3JJUNvBaqHc2xNVmj2A5Narf/WJMdSLcqi
Gkz2a/Pn/AuRWau9Muaa+mROMzsfzTkm4OVwsBtHiAx2RUIMqCNbyx7iCHJoNfyJNbb6tuYpBk3d
nwgewl5on27fST4KCByMqI4IzQ6+RvWVW6OXP7WkSjHtb7Ld2rBzpEaMEPcLwr2/R3hFFvrlyyXH
qbgGd3oyKPoqvpq3ciSUMNFq0mi1D5Q1UC02yjD+dkMaNc6G/+julxRBARMx5jv5hbbSYLYQqduQ
a/NxIDF+TOP5mYvxt/Wwbk8iWJEtvPl+NGfdvpSO+ZgZZ+Qa8wVPVx48hMK/9peZHce9kQSvVw1u
yL3Ao+lNs7TU5SqUYxZaBlDeNjM/4rdo44mL6BajGmhmLYo1mqm62QjqE2N9kCtZ88rFlkK/H3rN
RAfl6mJhs7yYTzeBM9ksPC8iTUQex7AVW/l4uDIn2NHKFoeICIpNNjg6OLfQZX3nrgig0T9BPIk2
MMupjk/GxfFfk/AU+5hYuu57624oy0B+QiaMGVNtE0BxLGwdat7WeD0mFZ2ZddUzf7dbMoGKr5pA
cgJCP+LCSd7Kd0wCgeSw5L+U3+UQqDYRWQxvRsrdzc/kO4iC8rB+sNFibiQIOgN9sntJlq5HUr4F
jfGUj3w/aIZJ4jDpVCoNKqskgBseRpTho0a7DVSEE/E2MOc+3zn+Z0Fr5QA2JAHU2wRkOUFKM4FF
oDXAxItLGmgihMATEyKeILAodbufj0uD/fFw1C1itWROo+mLL7hX+M49ZN3kvJ+bq7nLWgkGg0+h
Ya16Z6trF1ZkFElb87K9PWq1ih35BstaX7MyZ1mBiXlXTdrofvpcUsMe7mWhRIVKT5DWHPisAaOm
/vR6ryTvCOmpXehceLjAcbN8SFKHSk6D2V0kDJox1hVV/YRo9LaQ1vlE9EIRwLDt8tgGoNIfZ2l7
tAx9luZ9dCW6YUjQ8UiICJBTLXWKOj2cmhUR+7kYlbS79XHnAHqwNLBZwg/FqLHrkQyE+AAuUl5B
MXI6WSwE4Z3HvWKicDxBo6bRJjmXgwaEJlp0DHx9i2AoLhV8Jfwfvsz/68vc3BXSIKdI0/heIOf3
nLjXaGkUS4WZvkzE8JHEpVdF0FHUvwGOgfMQEADV1+CpOMEfRHYXl1tTnJOUOCmnP+mrlPjPteTO
80EaCJNos2ZZnzPZGftEeowS5N3XJeHmr+RZeCNB/h4n4IooUoUnrnP9Gm+PPJ3rD7r528IjjdO2
zFYrEH2JKwn0HLojdGnRYa6crt+NiqRYrT6XZ/Mui0/rqk0oLnEUOziHijHJDXYv4wOi2E97OZWH
WmZ6AZ1lAKT4pgrm2UJT7NIyv0x66Enj1iWcR75QmHH+QI3PQzvol9rzKDTtjB6JW2Vd/Hg5uFfx
eFWgipN9ksGU4ipf3EUJxhYcE//zwq4aqMX1EEJNIeJ+c0IqVNalKmNXE4WAWGFGp+rIjCKT675n
RlSaquBWSDEj44CrMwBT7mrg5i56xdGds9uPQh3IzaQ4ke63bWS7ZcytNInVIuJ+8aJXdMTh/VDn
hCLz3Uwk+Tv42mN+6giFbBKvfdlqgC7iFUeAOdH1VRvkLqHH0lUFPrMHEjfF0QA9z3ih0Mk/UoW4
Y5cGljpnAgHggKCqbu3Qpw/nrUvy8iwtA4iciu3TqYLBZYdAoRvrExDbFeOqpqln5tAATvrjRZyS
Ld4KWagxpitgy6exaNFnvL4ZutHh5oIe/F50tPn22NkLYicKoVRujRZ0eePU3mvRzaBYhrzQ2pT7
o7YYUjtefYg5s19ZYEaJFEkzmt335FoIVhE8NlnhZgxd+5PhPGwGn7q4nRldkrJKSgjNjHRqFiBk
u9bi6eSeD1Xd5YI4SAXfhNhUU7FKjFlwScda1KgMa6IQ1JB3GlReE6jzI7oySBRc4w+UI299YFOL
+7aumQzYBT3Qzqg0Tggfdo/53rI/IfqFcnxkmvrNL/e8MgJVmf5nEpTtgchZSi4xTL37aCSqf6Z9
EJA820hbXMMxqGPPYfU3PM3Zd3XNrnA+yHslVJG9taNrb+ftWxk2WR8GinU6i6e2CO8j+wecro0/
rdQj+mzNkbdEY4G+B6njNhTMp3ieCtfu6+VkE8ffbT9fxeB6JTyirpOkWPmMwxNtThaguNL/rUjS
XzwNv8iNgwUyKFIDvmhPTio1L2iAdTevwNvqrV12o6puJ5jl4bNFhTyw7gBwpCnHjmu1U7nQeBE/
VOm9bC+8PDuwuGdCg7FlrKyZXg79yae4DHuoqFXikWQUem8/pIwc9O1u89oIrXLyuu50+gLFjXOZ
SZ1hWkU4fcnQ7XuL/8IFEKVljjylmCPCNMPzIW4xK1SJuSyRmb98lo0WRAKAAnxzqe4Qx743VxiJ
ElNY6GMiUcCtHedYrf2E0DQPUwe5MFPo5z31rqInqk8zI0KWKNVpNOgfrpuHXwbRtP+6XjPAxhA5
KKbir00AkVrMrdxOXW7NINd8PoFfHYQcI9QR0kc/WyPXZ4Cmn23GFXZ3QRttFRX2ASAQvQxjGQBl
TMb83GKX3rJsKY+HA2RcPxiqppwcNxcWq0om6jUOFppQx3ziyzjpLxohGYh+VCa0GCBPzgv6yamQ
nNFWJ/Zdp9X+z3Y3Fbcc4nJka4wH1mwMBAHZNDT0Uc90l3ONqPhXtPZhh04lOW3a2/K/eOJKf7JJ
gKhzVP7/uqTg7lWjDHHKhYTOGOJ6tSqpIiWSARI3pkO/8IAnaBjgWOcdNTKexaqFlFzDBYwqeBQ/
YBM3tozutpUwFoVDPlJC48S5BgC8RfRqNw2VEYxT/qR7ZRmneCjCRJ6gqVpMFrIt882Q6DxlYy5r
jTI8HCDnX57M74sDvqx8s9M4XUPKHH/IDe0O3uEcReO8hda+1Rf7NELPGbPJ1EQuzMIY+mfR7j9c
QdhhXCHCuFPRS5LGHKJaU4eUgd2UHRE4ZSZ+5riOq8i7/HChgBjr12KBzlGFpUrXQl/n5IM2zd5V
xqoXaEZ/TNsmhUhBlpfquLQpn9dK5pVWjObi46c+nSZt2RLJvJi5m2MTBFvxJMpFTUu+bRudPB6L
5u3ERtD0sv36c8ZJjUx0iEeJKPRDyOnNV3JSBmhfWjma/TgYyF245xuBh+p8n2jmm+WpbyKbZndH
B+CGe+wjOsltTcaYKvz1arxAuqfTJVGDUz9JWyhU/eGqrLMW7uX9LJigbrypN2AqVjT5ofScAHYh
NPkVPG0IgzRJRg67HCOuSmHcBqC7Ib4QbJ74ECTsfeiYeB+8jjiT6ivQD6yEkEfN123rCt6RNDCK
9IWTtqrBOsnVzokgnNFnSqEqzNy258RlIXGR4t/GURKP640/kfiR5wbSDZr+m4wnX9kQcPu7iLkh
iWjjuu/AC0O7xLfJFkmqcKYtGfWfYAlAjVL9JEeiFXYYH+QLD3lbiqAKsFmLkYDCJPXKNaZujwTH
CtrCsYwpsUokNnwhLgflcKGEe32npcnqCyBsMCfBl2KpTRpoy/d2L5G9sFH3RRE0rJDsUFCjTPEK
ai0NQBBEi/K/BUEWN68xsnZAGL5uxtUT5ZgZ8TDn6PZsuKEfVgKRDzPi1ZkVBSntjzFHGEahT7Up
SC+VIEUjVkVFoRD4i6PFMBPVissNXbUFd7r9sN9ykHSbui3CG5AeyXpfCKUTlBVPio9MknbkDtG8
UEdfM/UA5S6YYnBD+hl5pS/OdIEQqi8D4YDi0A2ByDh71IeZnBv8P5DekmRil4QAbtXp7d4WzzEA
dWcOR5Dvojq8uWW1xlJwos1w9zRBRnMvuHONCiU2Z3R40pJ8dwcIkixyzXHQqhrEn57uD8TypVIS
YiAYTf64Nm4CM9ifwicTOGdvi345/2XFuyNYMhL5TrhuH/CUdCa1pnS4yzH0wVVpv1pfbVrYI3qm
3/TfHMiUa0vBTOuUFd8s5Jz+7wPuMyhPHrfggjiNEoonGLRI2C7iPetsbjD3m5v5py64aO8UNHhQ
ljmXKryBWUb/PuYcuOPiXt3CfzdmTKrP19B/3jRbYrO2U/+iEiKqLS7CPsSDPWOyAKoF/9KxHGD0
bsH4ccQ96H8bC4U003gMMzzTASE6udapPhgeMt1CxATB9Qi9INj4Qu1hQ/EbHVKnIOrPCFcRAmDh
1rCu6n/GoUcJIqZ2rnXs5fQCBuArlwMNx8B23NmGOfPQqgiSOdjEMJuIuTXUUzx6OT+AWqEyM7qz
7DAtACiRR62U13FR3Fv3yvxe5AUOlfAuM4rkDdmpIZHkAw5qExIxIY8hrCaYfu1xkC6qywQNxjNZ
Idl01DALTtoXPqGDCCyqhDtIshzKJ6jqfTgGNjF5QJr6koT6q1meJFVrkp6nxGKNCSJvZvAHWNDY
MnhvwAxHyE702ILzKj90m9rmT4zoc5NbeVuei2ltz/TiTcmxyH1khsNhogs0n4gtPPbD7kWOu8Uz
q/jZ1FfcUOKCPTyMjOjSM+MPMQom3O95dAMU7C4W7rtH8ALqMtpEP3AuH1/byJylague+pos48rp
xVx1CIdOds9ZTTrApwqByaXockBXjqQZ6MqWdTSKXG14AntHApHx/5j5fDdQCNNlE9z0bZmT+1s8
2vMTtwbrOuHN6KJBuJrRUErrxRqPrRefVY0dZOytW+031UnNVK3XdKQnvJ7LYB5Vv+LK+FRaco2B
5g8wDVZH4U+yhdXb2oiI4MDokRyNgM/CaoHxiBvCtNqjVplqpHhsNHX0rmeUK1fnt7M6YNuGsnn2
E6xHcft6HoAEru5RHhia6C4Z8ceI10juvUCOsgJS
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity FIFO_SC_HS_Top is
port(
  Data :  in std_logic_vector(7 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(7 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end FIFO_SC_HS_Top;
architecture beh of FIFO_SC_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo_sc_hs.FIFO_SC_HS_Top\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  GND_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(7 downto 0);
  Full: out std_logic;
  Empty: out std_logic;
  Q : out std_logic_vector(7 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.FIFO_SC_HS_Top\
port map(
  Clk => Clk,
  Reset => Reset,
  VCC_0 => VCC_0,
  GND_0 => GND_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(7 downto 0) => Data(7 downto 0),
  Full => NN_0,
  Empty => NN,
  Q(7 downto 0) => Q(7 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
