--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Wed Nov 08 20:18:52 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_basic_kernal is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_basic_kernal;

architecture Behavioral of Gowin_pROM_basic_kernal is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"39556CEAE29F59569B269A2452FA5E4BE8F66139EE05AF5456BC890C64A7CF5E",
            INIT_RAM_01 => X"D132A248E13A3129494AAD2D998C21E85714F9C1E8E9692B548A459F57B2C649",
            INIT_RAM_02 => X"4ECB54AA652BEA68E691EB2745B23A94DE4F169CE689BCCC5268CC4B3A39E52F",
            INIT_RAM_03 => X"9052C5215529839D1804AF77F46F80E2564448FEA910110154EABA6A9A8A74CB",
            INIT_RAM_04 => X"EE0E42A2A949E2EBEDEBFC2B6D820A248C990960364CB67DA20B800D4190C001",
            INIT_RAM_05 => X"8D03A62DB311F9631102291B3A1641C608154370589D09226498C87519EB3250",
            INIT_RAM_06 => X"FC773A00F32175B9A191896B07AF8A800919999E90AEBD98B30664796719EE10",
            INIT_RAM_07 => X"265C93290A5694490C121B21446A4A9B5D992C9C9361A996C1410A6ABA49B31C",
            INIT_RAM_08 => X"A4C96450B479ABE231496BB681364BDA0A44339D41455866609161A3C12AE0E4",
            INIT_RAM_09 => X"05414448211ED3204232935943B1EA809BFD00396159A612B5AED4A422721010",
            INIT_RAM_0A => X"503C4879AD9D16D96287313A58244D306B5A293072904DB046A949883B842122",
            INIT_RAM_0B => X"C6A58461D7BB32D4A272498A4B4A4988E24E4A2E19916E6CDC56C8008C102C2F",
            INIT_RAM_0C => X"341BB151A2249685044A52673A6514A44994ECE68AA51B5C518428239345A4A6",
            INIT_RAM_0D => X"81A227577165DFBBB2D5B008112A1229469F6B7F71511BD22908A1A812B1555A",
            INIT_RAM_0E => X"25C1A65ED7E89893332636506E594B63D596592D320CB2D1840CDA3183710142",
            INIT_RAM_0F => X"47FDD0B07F4502059940484918081C44254530890408842022994A7A8EA84A52",
            INIT_RAM_10 => X"79861869422F51B3C4D25A444B2C4040862229444278CC81318B511AED37EB7F",
            INIT_RAM_11 => X"FABA85A320CA8573CE89380947B1A17B6D9D786992B4999C1CAA935C8DD8BCB2",
            INIT_RAM_12 => X"3C877C3A73D452A13024EC86999301B1C1A5F0082CE4C8139B1A6CA166759429",
            INIT_RAM_13 => X"45ED2156816C92B2513290260130AF416A98910006F9C676B202B92B050692B0",
            INIT_RAM_14 => X"8DA02840FAEA80124888F49933526438110198C44444652594674A5C03326996",
            INIT_RAM_15 => X"0AFE6588120514853612A17084F4A88922E27E6D6127F69933321986C3019D90",
            INIT_RAM_16 => X"021661E98201E5441110A6703C1A0833320060484A962D9171715693D5DC79C5",
            INIT_RAM_17 => X"7CC5A20909224A94050A8A091084210A401E418577881688D7CD6010A025010E",
            INIT_RAM_18 => X"4E8A41410069DE977A57455495810384187048187AE856350D22C46991316C95",
            INIT_RAM_19 => X"3AF109405A9087661008A88483050412810103BFBBFBAE88823FB044715FD5FD",
            INIT_RAM_1A => X"00A5020222D3AB4235BD2BAAD2B490110AFEAFE8B582B4AD3BAA50B852AC4EB5",
            INIT_RAM_1B => X"50E5D394E422080D2AB4AD257AFAA3100715FD5FC0110C3450050184BCA04906",
            INIT_RAM_1C => X"E901BA3F4888711450C733A11AC4D74A352B4282480B3AD354CCDC34588A2116",
            INIT_RAM_1D => X"8194A5E0D321332C9CCC520890CA2D402441122E05021CD5920223133918CAC8",
            INIT_RAM_1E => X"B5D925FE481A44E003A9927941B80035FED7EC264334252CE5C910200AC14F8B",
            INIT_RAM_1F => X"0A5161138C2DE03C9D30C06124844C0564B0000000001C1D8FC1D0C941009AB2",
            INIT_RAM_20 => X"13096BA9B1B21070D6B45291891042146B18302FC60D0E19354C4B2EE6B604E9",
            INIT_RAM_21 => X"9004801011956D289612490EABC932CE26C4856A651D3504D5CBD04102184405",
            INIT_RAM_22 => X"ED9884E74C21586012C472218ECA8815A060C21D0A0130022B000428B32480A0",
            INIT_RAM_23 => X"A69D7C74393B9C6A98948980432024036063840D61E3071F5201B29D36E44EEF",
            INIT_RAM_24 => X"42D0A58967040BD6DD9191CE6B00F057C01B8D3C25715388395B860C1608B0A0",
            INIT_RAM_25 => X"E1388C2849A2B0083224E6D790543089C1A2C2063E0944975A52D3B76C448900",
            INIT_RAM_26 => X"D0497ADBA8051A277C80010800925D131C3E5056B024012BFA421D2C590049C8",
            INIT_RAM_27 => X"A87A615A94F0803103096201492E5E2A2CED36D845B015086622AE5CA1950440",
            INIT_RAM_28 => X"789966AD2800302015E005680441031424910C61143D1A18B20D300CED36D858",
            INIT_RAM_29 => X"13F96FA84DDA6781052D95A8AC144CB202002B05960DF78687988AC2224B645A",
            INIT_RAM_2A => X"3703014E408944366780D82BFA918680D7E2380E143C35AADA985DF6E0D03409",
            INIT_RAM_2B => X"0EF4A5CD1C479F5B877812E68E23CFAC371BF2285330DB1C31020A8081421662",
            INIT_RAM_2C => X"00002B5528040C0001FE96B9724710EEFE0DE73641CCC99E5DF113A8F746D6B7",
            INIT_RAM_2D => X"DD681A21048401AF46032085B7B4ABD04A150B744A522428482B42B689009200",
            INIT_RAM_2E => X"282B3E858F6F7EE891005AAD5EAB57A1100A1690B7482846C14B69EF96E04826",
            INIT_RAM_2F => X"56F7F7D3B20F80490D15E84A55906E5CA047D02820CF2D55457F220A4DB4CF20",
            INIT_RAM_30 => X"1DCE2B5218255F25F138500A84CCC101042B3991652961499911189C5014C890",
            INIT_RAM_31 => X"06454474B61068DE5D46300A254A2671316076C6BD84DA24C899D78DB555EB70",
            INIT_RAM_32 => X"D8002166F62B0885CC854325A609A1A9703306AF4ED6C0C21E1A923063B5829B",
            INIT_RAM_33 => X"B0F139E2A463A39330F6C14C548C56EB4635EED1402DA1A6A912B6B587028DB6",
            INIT_RAM_34 => X"ACBCD71A055BCEDD4AAF4AF09C6A3246672A60E0714C60530012F5BDB44FBE09",
            INIT_RAM_35 => X"BCBD31F51A384985ABC1A01820C21524620F115FD115B019EAB4868810442424",
            INIT_RAM_36 => X"58C5E1224C112141B20D7D0406D5898F2223E50A604CFC6A4845B22DE61B8AD2",
            INIT_RAM_37 => X"B37BDC4F67070A40FB204B78488DB7B1437406F3B766C3439D50211311196596",
            INIT_RAM_38 => X"0F18B136E478441A4FB7FB003B0C8F490F189256E0C5756810421F4262ABA77C",
            INIT_RAM_39 => X"000E95B8470CE50744F22024B0A0E5D7DD7E024F7242F4DA52DC89B002C61158",
            INIT_RAM_3A => X"1203228C84947071569D22AC00B654305A9974296B8B9004768694280A243AF3",
            INIT_RAM_3B => X"A75FEF11822D95926B066007439F4509B2316D81849A41E51405913B43738133",
            INIT_RAM_3C => X"3698090903D4DDEDF284DA6010A802019180201273A2A53C1E6064503102367C",
            INIT_RAM_3D => X"171A7C9C2FF7B80C8EE94F7AA8A540043F3FD1440A49D39BC1914BDB890549F8",
            INIT_RAM_3E => X"3A5366230419C1700EE03915618B799305604D8C050DF040208041065701B2A1",
            INIT_RAM_3F => X"8624CA4886124924C169364905B09A6D074BF1DC649340B16922B2AB409E9DC4"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"9A2AA43A9C6ED6B6040A201E87D67BD0EAE23BA5BA02D0ADF704544440E48ABE",
            INIT_RAM_01 => X"0813108D519459864C321891980A45C5644978CEE7B2E75D170BC94B669A8EAA",
            INIT_RAM_02 => X"06C0E01E66A88050434B50C423D1409930C76C204018DC4588BC4434941010B6",
            INIT_RAM_03 => X"2AB902108752892A401991290A80049CA188F06EFAABEBFFEA444125734C89CD",
            INIT_RAM_04 => X"502295C13A28495009045068282F2AC686A52D183489A25ADE222041AB0A8056",
            INIT_RAM_05 => X"41E1228428249040243A000022A2055239960809170A31408510504144241014",
            INIT_RAM_06 => X"AAB4002026615014049503222515040E344141160D012900A64404414C32B141",
            INIT_RAM_07 => X"00D01A29D4A114AA20D40051250306AAAA4301090B074C00D21218CAAB60E610",
            INIT_RAM_08 => X"429204498EA1045661711002C00092D2924082A15761405103A044008308A504",
            INIT_RAM_09 => X"883A1016290001280905A841310A107E0454A909608034108068022804D81ADD",
            INIT_RAM_0A => X"1088885A2C11C2D1085512281206C1A60000600C40020401142825485895A848",
            INIT_RAM_0B => X"9495504AC511A6A5365978CB442578C8B2A3024A411008405490D11CAD954303",
            INIT_RAM_0C => X"160AA14902842508D21014455220A41600A05544600572501C000B32A8460246",
            INIT_RAM_0D => X"90205A9150A4004A800D847ED628082019D0940504114438106B3428049D30F1",
            INIT_RAM_0E => X"002DA24484288C8154454D5A2A494830A80482A112412011383406020117DED6",
            INIT_RAM_0F => X"42285080B18993204A2C4AE01A2904E4A0412420450214002044821100040B54",
            INIT_RAM_10 => X"4504E0081A908080A252C85AC90108030559BA05D2A4011C1664050554254221",
            INIT_RAM_11 => X"040148104010A4001048080004610252490A4040802541101488885101002824",
            INIT_RAM_12 => X"A0482910AA09B00C812200E9950400E13D490C01A8846B713255080233283500",
            INIT_RAM_13 => X"89414830824835820DA2C8E2034B022D0982568B8810A40460F506B4932104AA",
            INIT_RAM_14 => X"0936300944092E185061202822544F8B0231080888884921224294942204D520",
            INIT_RAM_15 => X"D48BB8C88AA265085280FA890C081131DA29292041D9522E46CA0CC42A4C1404",
            INIT_RAM_16 => X"4400C15102CD45442621A81380044B26202C53060B0408B00A0E064682A10287",
            INIT_RAM_17 => X"016992E4080023C9F36AC11094C830BB6400100C014274D20168451D41802404",
            INIT_RAM_18 => X"90002AEFD82A0522400A10504400C151020ECA01155450083905C0EC00300005",
            INIT_RAM_19 => X"40894980421BA73E005F56404011440ADDCCC90411555515F98285EA8AAA8000",
            INIT_RAM_1A => X"0095B42120A5280004024554A108A52BF554000055B528420146D40440800624",
            INIT_RAM_1B => X"A10AA52105A90C82452842290055270FE32AA800157AC08100151433802A6DB0",
            INIT_RAM_1C => X"2A6014A02508002B2010C14840A80240A0401410035081A6242B0094C121A241",
            INIT_RAM_1D => X"209209141903CCA0EF58843340149A80120CD208F478A15621026228A905488C",
            INIT_RAM_1E => X"0AAA380181708088096129544151A85AB44081042A455A5A88280E9D48A90140",
            INIT_RAM_1F => X"0A0940266517FB162A8A9091A48854310681FFFFFFF80D1D9FE1D0D051C00020",
            INIT_RAM_20 => X"910D00431E4A2818912825178921030500448E08D1084B42204444401084240A",
            INIT_RAM_21 => X"CB0648360301622932CB54D492CD15466A8728025219AC06B190C845805865DD",
            INIT_RAM_22 => X"85B607BC8C528C48F465522A951010A5006E0289796D8D9B083984DD21210436",
            INIT_RAM_23 => X"494828D92288D220380454ECEB00AC5A203F19CAC07706ABD20882AC1024BA95",
            INIT_RAM_24 => X"A33004025A10122A8023118608E6A934DC0868AA2C5F63CC0032C408DC0CE0E3",
            INIT_RAM_25 => X"2AC64A68F12C583268E5C30A429108210300BA2A4A80104025A989628058B821",
            INIT_RAM_26 => X"8183002017D46AD5468218DBB2588022A8A35748113210AE8A128A81C1604800",
            INIT_RAM_27 => X"A80224448AA0B020E0C01A060921555A4B04240241A48D3A5400225403103876",
            INIT_RAM_28 => X"27D20333A1C45B8D455B514786EA3050D48C2B4D008820502EE3039B05240200",
            INIT_RAM_29 => X"290044440A08121A988AA68008A0A901BD44586024F00080542810000C402000",
            INIT_RAM_2A => X"045AA112C04B05484028011500888810311000410BEA587E010C0A8524250141",
            INIT_RAM_2B => X"AB21C79254E8CD83559C63C92A7466C03C2C4D1C204B140B6A7AD0858BD48000",
            INIT_RAM_2C => X"0000D16636040C0001B6FAB9ED9D3ABAFED25042300510AF1651BC94DB115B06",
            INIT_RAM_2D => X"9006000405248804211201280420410F9A8340035294A84CDB000680D1A00000",
            INIT_RAM_2E => X"A08080A840085420025A000008000200D10480240026122802501908A04693D0",
            INIT_RAM_2F => X"0040000902006480004C20BA44014880140006A644005254240028490801005D",
            INIT_RAM_30 => X"2825E4820E7665798B0A9C86AEA0032B6C6502540313528220A0822884154045",
            INIT_RAM_31 => X"802020207018501200C01AF182300229060600B1541F482808D00316CA9AB130",
            INIT_RAM_32 => X"200DB61090008880423111454E29A2240258062A5696D150408655B155A5B000",
            INIT_RAM_33 => X"20B000041505905280A029532828106A156A010753AD241A855809620858126D",
            INIT_RAM_34 => X"A8048A3632C81404CA8B5050E7CB20CD012821E071065811BA00420A20454528",
            INIT_RAM_35 => X"822D5A0368A14D04A2442C3300884021555584141AA107A52A14328EE408299D",
            INIT_RAM_36 => X"814500C1820012D00D68823368440C502B583C026A2040810835010003001692",
            INIT_RAM_37 => X"40001081017192F70806E21BEDCC050A1AA2A084204495728959218141004804",
            INIT_RAM_38 => X"A86004909916D60329480240281103540B2E0490460022955A1069E000110256",
            INIT_RAM_39 => X"222C963175C0114A38C2D820000422020A000A0200C281021001814490001002",
            INIT_RAM_3A => X"89E8C0A15821252A000D010766A30254902403020051278A54EA27526834C862",
            INIT_RAM_3B => X"1577FCF00204404050145E12CD80B400134041726510080A1810901248058020",
            INIT_RAM_3C => X"3009882CCA2001045244C0278402654403340AB808406909439752D012582026",
            INIT_RAM_3D => X"1D840402C44A1396D492001552188ABC0202245C89100F65EEFE09428C231924",
            INIT_RAM_3E => X"A354000200800A408110002028D9424053590409148021435D64F3C80003050C",
            INIT_RAM_3F => X"9DC21A69205A69A6130090D34884402DC810060484D02202A706116255310504"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"2BA7973B6B976ADFEAE9A5B7DCBE5000FBBF547194BA1479505510145C578041",
            INIT_RAM_01 => X"EB77D69FA3A7FBB75DBAD695DEE9F816BB6B11F82A46DDDA6FA1E3FDB4653D86",
            INIT_RAM_02 => X"6CE76ADF764529A57A83140ED024FD3F9EDFDD69795BADD5718DD56BA75ED6B0",
            INIT_RAM_03 => X"A02800915229029D2C008B14A44080226A4848B151501101144015B4F5DFFB9C",
            INIT_RAM_04 => X"AE0C83441161E3DFE9EBB1460B260161822814121404932D6081AC0561806349",
            INIT_RAM_05 => X"08A0062D308400A121091A88AB862547967C03404A04080A02ED9048FAB7E10E",
            INIT_RAM_06 => X"EE14998EE22459F5E4044200A36C8E00312BFEBE8D9E1008A214C0594E699519",
            INIT_RAM_07 => X"44405F028A4208003E0A8132410015585B9B4484880120924242094B29B9E210",
            INIT_RAM_08 => X"A24925E620688A76D9286E80E022490394405D5F993A01ABF158428C47402C32",
            INIT_RAM_09 => X"64A13A56A44631404337850467FFEFA5C3F5E1407585372004EA060120FA9908",
            INIT_RAM_0A => X"308A0848950910036BD142020082D59A00004508EBA0FDF1F32B8F10177828A2",
            INIT_RAM_0B => X"5250C4A8D21C863013293AC1C1013AC0117D5726ABD4295A0944440D80442502",
            INIT_RAM_0C => X"B3A9018ED800862102FA0BBAACA03944C05564762130A10D115205DD551A9168",
            INIT_RAM_0D => X"51A026E745D19E0080C801147D035B0200E94A5713012E40721C82809935D770",
            INIT_RAM_0E => X"5269C991B5A00B80B00144222A828309FDB2491C422496E0943DBC00016289D2",
            INIT_RAM_0F => X"25F749BAE709C30D9B68401FFA809BEE341589116F2E5E82B25FF866066A5C20",
            INIT_RAM_10 => X"59CEFA10580FC123AA00021E500F0201BC2028A5C2E604F9EAEF0A02D90BB95D",
            INIT_RAM_11 => X"73888D8360DF4840DEC1E8050F138472490B58E50A22ABBD45082F4408442CA6",
            INIT_RAM_12 => X"AD851872634CA0945804665551000C20A16172446A559E931A57681977EDB240",
            INIT_RAM_13 => X"8D8FE135C12CB1B04887304238B8E56C630882C006319656908639174C82BBA2",
            INIT_RAM_14 => X"35363CF8AABC8E3E04A17201BA4AEE15CBE118C888882541B4658C4A422471B6",
            INIT_RAM_15 => X"8A77D5CE91AC0001061951600050A000BC65514D72BED6B5075F35C66B07E8C2",
            INIT_RAM_16 => X"A0304199C958A0D8000117F33C10052222C8FA2CDEA42DA3762A5A5D45ECBBC2",
            INIT_RAM_17 => X"0DFDA15610446174AAAC873101202190C01A418D674004DA07784B88A1170084",
            INIT_RAM_18 => X"DA40EFBA8821428D1E9E00585424617A4A26B140BFDA701618018843B2336FF9",
            INIT_RAM_19 => X"48921100B581281C0235546440AABAF788D9CB3DF6CB3D9F519290BE8D557FFD",
            INIT_RAM_1A => X"82958019B2B7912A949427F84632542BFBEEEBA008D2118C2BE2222C40001204",
            INIT_RAM_1B => X"F221B08C72C58B1426118C95EEBBF990219557FFC52FC2107DE28A4294491181",
            INIT_RAM_1C => X"A181EA7D07B012153110130C0D8CE61C182427447B3AF89118098914890B4216",
            INIT_RAM_1D => X"00E21D460F40AB007BF5C01863065FF32E019B8CC4683D9F713068028815022E",
            INIT_RAM_1E => X"00002084C160809AA1352B50E1140A3973CF8C1422483C0A01905AB1120A470A",
            INIT_RAM_1F => X"30114007C2EB9F503B90C080B10B5A22208C000000061D0C0FC3C0D151000021",
            INIT_RAM_20 => X"B0C122E6EBBA00400E10C24B0A20CB24A228541C4A49082830560F156007903B",
            INIT_RAM_21 => X"A8344192818244083CD517C3EAC650C6A6DAE48A1E8CDB336CD0D06596184F0B",
            INIT_RAM_22 => X"84AB84846649C04882025820CC9898019B2CB20EB325140A0110A51C3161803A",
            INIT_RAM_23 => X"1B151026D0F0240F18040146114F4111300372C4771BC9E49C0080245070C8F6",
            INIT_RAM_24 => X"3A0904C40C87F9C40401106BE304035F8013A60021E7DC751B4B51358835E373",
            INIT_RAM_25 => X"A776038C7DA3F83B3234F644F0E2F82508817D021800201F88E26233243E7808",
            INIT_RAM_26 => X"459038C897C46C253A0011C1E21833022C3B030C9390B83EC44015198E91401C",
            INIT_RAM_27 => X"A60EAC9508AE3A18CBC11D16642B061CE18580012164AE3745004B9A818FB436",
            INIT_RAM_28 => X"679B6C3BF8C2330D04C34121D3E9F900DE0FA3CE802C8B0C1EE393D18480016A",
            INIT_RAM_29 => X"122D61FA42286431C4199C80FE980DB77314316DB6F451820C8A0F600E4582AD",
            INIT_RAM_2A => X"444699696A880236152168B660AD4601D3320A028DB1783DEB38C15012C10221",
            INIT_RAM_2B => X"1B92734315B5283E0DC339A18ADA94EF407394064319C35B38EA6F66688E7141",
            INIT_RAM_2C => X"00006DF84606080001BEF79DD0CD6DCBFFE4D012398901A87736F8A5B4A1C87C",
            INIT_RAM_2D => X"B52E1A2D612489AD66188503FE7AE950D8970B7310841D4A9B296526788D4800",
            INIT_RAM_2E => X"AEB9EF8387FCF60F31205AA55AA956A3C32E16F0B70F1A52CA47FB9C2675C834",
            INIT_RAM_2F => X"5A97D75E971DE6214F0DCA7CF1C4607C1605F69F00E53E09617BC39F9CBCA739",
            INIT_RAM_30 => X"4F4E0F7B5A360A25BF18C02C8E8AA61A24CB11D16B1F41E08208809A4EB94010",
            INIT_RAM_31 => X"060000203F5D0A9644A5260A055812125345742BA897C3AE40915DBFC9DA75E0",
            INIT_RAM_32 => X"43290B34B7390496251D75102205E50D383E27238AA2F2C74C09C13C12A89A9A",
            INIT_RAM_33 => X"82F930729622F16411A02C0C3E2A86595015A25683C5448E1C22169483120D10",
            INIT_RAM_34 => X"48B7FD1C07998A4CD3828A27510B40AC55CCA07C8A7850A3511FDC94F0EB1BED",
            INIT_RAM_35 => X"D00A2555E4116816AB55BDB3A0931672A0380015D601203DA0F7261CEE089429",
            INIT_RAM_36 => X"21E522A54452DB02D56911232541994322004D0A58684E475025354DED11CE54",
            INIT_RAM_37 => X"BB5A964A72810067538042BC4881B1A0F196A6358F26B227A28C41011984DB69",
            INIT_RAM_38 => X"890855B25437F0096DEF6801ABD5E84B682BF780AC2F33154E7033E0129B8C31",
            INIT_RAM_39 => X"0220101661807EA736706AC6120DB579DF13C12708CE90260034009190C2402A",
            INIT_RAM_3A => X"3001820708C41420040D05670011CD484E19C6789601000D72CC367880E6F581",
            INIT_RAM_3B => X"300A0398E0459CCF78F278825AB746C88A0D2DE95609E0C356804F0940518793",
            INIT_RAM_3C => X"A69193099BFC44FBB4A89A47E16002B6DB5B2A7AF8A6D6BBB16804850106723B",
            INIT_RAM_3D => X"6FF9EA786CD6B55B4FFF2FF000C4C488020210294000FD71043C0428B50440F8",
            INIT_RAM_3E => X"3A844AC191156D840E79319479D351D3475CC989890FE01092632CC657A19095",
            INIT_RAM_3F => X"A82DF593FFED92D9B7DFFFB5FFEDBEDAFC3F3B086360C0A18F2CDB8C9010C5CC"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1850069A48044194430C305485B37BEF1151D13C94FCC596F803FEBAE8EB2444",
            INIT_RAM_01 => X"B01360CD0188519A4CD26335919412102C49926820039D5F07515041A5246CC3",
            INIT_RAM_02 => X"ACC54067631162091E53AA03040050015A4586A11C08886904C868A288475319",
            INIT_RAM_03 => X"38D55A2A2C46394A82570C18C684FC86F0CC40F0510551154040053A39008D84",
            INIT_RAM_04 => X"55884428409359715B011009628A22818E186C68E70907043C8003D20A740844",
            INIT_RAM_05 => X"CF45EA34E338DE4239F60B133A184D8623C853604050271208510ACF50360A95",
            INIT_RAM_06 => X"B8673A802ECC50181985C86B05D744FDCB0150449534EB592ED529474452E711",
            INIT_RAM_07 => X"7788CD0715AD79822895AEDB606A5D030CDB3B5B717FC5048393DAFA3090AE91",
            INIT_RAM_08 => X"5CB6DF26BAB924D0A2571176717DB64D0CC6AAA894160F5556AA4049B722F9D3",
            INIT_RAM_09 => X"EC130048AB5181634F6D9A5400000012181803783819D3A2B064D68655050191",
            INIT_RAM_0A => X"531EF973098114D06AD6751052D1D8AC463020144003811510400FB01C0D226C",
            INIT_RAM_0B => X"81E047C1919E26F483191B40C9411B4042AB5983D1100D7E878785900D41CA6D",
            INIT_RAM_0C => X"57B0828058AC6D6B1CBA55415CC5297051AB9890D8215A0111102A0AAA403C0E",
            INIT_RAM_0D => X"B3839364357114D11A989E288902BA035B718C663F1250F08DE6152010311468",
            INIT_RAM_0E => X"7FED4489CE2A322352776E32EF8282588B6DB4EC263249364327F499A2551744",
            INIT_RAM_0F => X"6A0851B839F97D727B6C43D0F020006E61450E6147883428A0900208C89F8624",
            INIT_RAM_10 => X"4104501320B09012C410C01470224043BE1C28AC1E3063A5400A4F1D710C46A1",
            INIT_RAM_11 => X"424CF24499B5EC3246C0080A84E441D6DB58C05A551D01100F2A9049E78D1BA9",
            INIT_RAM_12 => X"A2706A5122305501044BAA80575DE9AF19190020C88106817690188022BB646A",
            INIT_RAM_13 => X"9B0F4072F6D373321C01A1A6681010804237701F84D681A9436100A032A8492C",
            INIT_RAM_14 => X"03E1CA0000060110C81029120AC050000001F8CBBBBA5BC56E9AB5B4ACD5916E",
            INIT_RAM_15 => X"010280880880CC4200A2001849A346600402868440142000320A020C82180401",
            INIT_RAM_16 => X"7853802450201C41CCC2803003A1D0EEE3A44902040C1BA48ED6A2A092A34280",
            INIT_RAM_17 => X"243C32803118120301540C058330830084E13E790181F058D19C86A01E817C20",
            INIT_RAM_18 => X"008E0000464008102043C4140980039006D0735B9466B2A8202240A24C04800C",
            INIT_RAM_19 => X"23C61A00001C466C06C000039640000180044186186186000087080034820820",
            INIT_RAM_1A => X"8009033BDCC1704E0D08CD118C6001940411555AE9F18C63140CE69D92265EB9",
            INIT_RAM_1B => X"2010C842006A030088421002910013CFE7E28A28A455542D905104D102E35917",
            INIT_RAM_1C => X"EB420140681845004AC675E1C5C203C10308001800A003C84C4E473040B06148",
            INIT_RAM_1D => X"81A0C1E09F681585F7FD9C77E0DDC8B77E791682A15A2B15EB1003BBB00DC0C0",
            INIT_RAM_1E => X"A67BE94FAD5CE6C20BC1F27E1FF988942870F0074BE069BCEF1B56A91A4B5CEB",
            INIT_RAM_1F => X"304D60417BB3518F0C0BD8F7898F542E449DFFFFFFFE3D0D1FE3E1C149C012B8",
            INIT_RAM_20 => X"434A080800041C70C8420801030D2038118600C081C56703654C80608B19A198",
            INIT_RAM_21 => X"F616808045964928884F0D4C638E230C889509A3740EDB9B6EED184112194312",
            INIT_RAM_22 => X"3B5C05CE7E68182090E270C38646A4393B48741E0321AB034220106433C5989A",
            INIT_RAM_23 => X"9B224686030124C9C8DCDD88C102C928701E7CE6B15DCA3454C1183D63211D44",
            INIT_RAM_24 => X"925DA01104232098A8A7B12A03E440179C1201100934289C3AB4C2A9150236B4",
            INIT_RAM_25 => X"CD3987C8354301C09611FE99226543CAC27A002EACB3D6BADE76D3BE28020148",
            INIT_RAM_26 => X"1C5A473368311427011FE2108482449733CC041624040103003EA22050129102",
            INIT_RAM_27 => X"804062991CFB9E83283F2C31124C0824208C49261841924466234C803E408D80",
            INIT_RAM_28 => X"78B6DBC3F054F02078201E08F010C2C52F96058665311141C004A4E08C492610",
            INIT_RAM_29 => X"06C55B5412224DE8D92E89AD5E8CDB6CC9D51A8B6D0984AC971AD56A628D446B",
            INIT_RAM_2A => X"370F18127AFB1C37324D6EB98CAD86BFE18120499892501892AC34010C9C4548",
            INIT_RAM_2B => X"0B97F7DCAA0041FA05CF7BEE5500201DD4CE7A7AD7198B5C919A6CA8C1CC6273",
            INIT_RAM_2C => X"AAAAC9800204840001B6F7BDF62B8999FE64F714DBDDCB3A173DD60ECDE983F4",
            INIT_RAM_2D => X"FDEEA6420DB69C2B7179A9A7FFD42BDF90816B4F5AD6886B936F67190862DAAA",
            INIT_RAM_2E => X"AF3BE8878FFFBC6E836B5AAD5EAB57AC8100D686B4E33254230FF3F5B0FF9B74",
            INIT_RAM_2F => X"56F7D97EA765266D6F59EA14E5D146F4B65D060336ED0205754B43DC5F3DAF8D",
            INIT_RAM_30 => X"AAE7A0F218238221FF38400C30CCE25248423AC1E73762B139B310ECBE898C9C",
            INIT_RAM_31 => X"2E4546708F8634CE11AE16FBAF5A146A3371824C453D54E0939DD795744C59C0",
            INIT_RAM_32 => X"DC562B7673C2A0300B991334DA40438C5AC7F9259222218F16B3C4082488887B",
            INIT_RAM_33 => X"A20E19B4214C74E18CFC485A6E8444980319CCE994C449362C44A719A668AD92",
            INIT_RAM_34 => X"481B88B43292D095102490842AC03E366648E504165CA3A1E25FFCB4FEEB9A43",
            INIT_RAM_35 => X"249244034E08191080552A1CEEE90578875A158E5537C7E12AB18688AE688D98",
            INIT_RAM_36 => X"6A69881020DADB1AD00CC4800145248D414184681AECF68B1941340D6B1AD204",
            INIT_RAM_37 => X"7F7BDEAB74828AC55BA6ABAFA55DB21B00CE2E37B30048071880471D51BFB6DB",
            INIT_RAM_38 => X"04F25C000A084284018C647C1A090410045281F268606648AA123F5230253FBF",
            INIT_RAM_39 => X"788B372C4718856AE8F66AAEDA45788CA04600CA7B12E3EA31E9A04523CB466E",
            INIT_RAM_3A => X"E3F3408D77A07053679D2D5C64841244C093B455B19BE79A448AE457CAE42F7E",
            INIT_RAM_3B => X"B75F7BE43AC93914536656A7C02231737A354558313289245025DC3253738632",
            INIT_RAM_3C => X"F490937912AA1069A4BDD243458274B6DBDA00800897024C04082D81F3487CEA",
            INIT_RAM_3D => X"51EB5AD62637ADBB4FFFEFFD51A7D32583030181124D4954046A1210830C10F0",
            INIT_RAM_3E => X"BE023600C39880BDFE7E1BA1F0127AC70774A908890FFFB8924124820238B32A",
            INIT_RAM_3F => X"EA0B2DB6CB6492DBF6FFFFB6DB7FF6DEFD7F795C51227FA009249B0984CF0DF1"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C44AA1259758B4690471C4C833E0FF7DEAAB8429FDEC44155B12051142451205",
            INIT_RAM_01 => X"03E407125A0422009004082040228445C0A26607D5E43E10B82623220B899134",
            INIT_RAM_02 => X"9022880010E48790015052C03AB08580E01A2B4C01033194ED71959104000006",
            INIT_RAM_03 => X"E357EF662CC6610AD06A4890851084101100B000401115445151110944805210",
            INIT_RAM_04 => X"11425832C48450401D0018A1009ACA80C228A40B0440A204204658654DA19624",
            INIT_RAM_05 => X"EC59B327446ED919B9102E6664C337242015C288608105A348004B6C05254A31",
            INIT_RAM_06 => X"21041059B320E153421229045514542C295405544000448DF32E93F1E402A79D",
            INIT_RAM_07 => X"2266602135B583C72914000A048A500008010909610410231B7B2854EC0CB37E",
            INIT_RAM_08 => X"58924050482D045A04D6D540010492420960AAA9358081554AAEC010210B0704",
            INIT_RAM_09 => X"455140646188436DA100A0894C554501710740810262300AC22112708E000093",
            INIT_RAM_0A => X"1ACB3D40607113426C5D8CC74014439039CE6A0D1590020A0C9E4C44380D3141",
            INIT_RAM_0B => X"0C836124CC910292224148CE000148CB22A902985133C84830180E09341210B3",
            INIT_RAM_0C => X"D22650302C24359C6049540141140C9484A2120846C54836900CAA00A0810802",
            INIT_RAM_0D => X"001202C99A24200CEA0080299594A82C54139CE39F1A007000A840444D883081",
            INIT_RAM_0E => X"00241B26846EC90949998850183B2800000002008A00003200200211D395307B",
            INIT_RAM_0F => X"6000C082AD44830001248840D99800684272B088890890CED42004002014484E",
            INIT_RAM_10 => X"E2340464A2000ECC93DA394007204358B4C0655A222112080040230046B00003",
            INIT_RAM_11 => X"4208C0300801BD0C2048182A240010DB6D8C610A544D51473044605203264AF0",
            INIT_RAM_12 => X"700A0C98B2B75E68A198BB0A998090304383840D1C36485997788CE628201188",
            INIT_RAM_13 => X"40401A11124014848522929364014AC886C42D240518C02930084248211D1471",
            INIT_RAM_14 => X"6B042100888A4A46A346894C45410000D41918044444481400025296311A0800",
            INIT_RAM_15 => X"21A800B9CED912B5BCE60400B6A54888119AA2BC8C011C6022A02AB04C85533C",
            INIT_RAM_16 => X"8230411330135336111180026AFA201111491256CA5A4000115192AA82982C00",
            INIT_RAM_17 => X"C66582A919320603155988CC148460124054810499790CC9114BC922112B0B7C",
            INIT_RAM_18 => X"8021100026444891226A886663424101A505667A004494C30CA08C4923324A0D",
            INIT_RAM_19 => X"4088B3C0D695E35C05155578288AAB22022235441041042004424E0118000002",
            INIT_RAM_1A => X"004C19D3618064374E010002108406C00000001C23318C6340068C8C902354A9",
            INIT_RAM_1B => X"04848210806049210084210300002A20124000000A8023D202086059826E6815",
            INIT_RAM_1C => X"1D8001800059018000CC2110A6911A22C58288A200C40080081826E762CA6594",
            INIT_RAM_1D => X"508921880B4C158831FEAE54D825003226A93313A3D9EB35289A14444D626911",
            INIT_RAM_1E => X"846C4108A2C138E6410986710012DD1C3870F0269316A889131A7668BABF554A",
            INIT_RAM_1F => X"11A940F1DAB0FFE5084490238B82260C9CA8000000021E1C0FC3C3C1D9400234",
            INIT_RAM_20 => X"4D83040000042810008410819E11642944D4A9A395094A530146D59541C93212",
            INIT_RAM_21 => X"C0060010C184C11892011024A6C40976B3C0200F008000200000C1C71830E521",
            INIT_RAM_22 => X"0B140508480A084804401940D524460C1240240C110180031000300CB03482B0",
            INIT_RAM_23 => X"92282366080A4A14616A3099C164902A20229DD76B397B7D9960402948321046",
            INIT_RAM_24 => X"22262628600A4802460900D4180A232000084B083120280410864400232AB436",
            INIT_RAM_25 => X"31613220027409CC36266C8800082C5C2D17AA32BB84E000000004004050A508",
            INIT_RAM_26 => X"852CF199BE834159D49826484C202246682124911821646ABB8548C5652064E9",
            INIT_RAM_27 => X"193BB92249A002E49687C214C93830C99C6336D8408364C84C9891350914264C",
            INIT_RAM_28 => X"228003FBF41962698B0262C015102F0C8000180103E064326BB90C2C6336D841",
            INIT_RAM_29 => X"207310006DD000482C7B449185424000A00B0F4000A8A2663D8918D933643321",
            INIT_RAM_2A => X"CCE2C48C061C808089B7209441A4000101088030800C07822448A2A6E801B104",
            INIT_RAM_2B => X"0BB3EC230B08CA1696DA44139796770A81A730858DA460483406003004211CC8",
            INIT_RAM_2C => X"CCCCB00000020C0001F7D7BB09CBCBBBFE0948A106B226485775E267DDDA7C2D",
            INIT_RAM_2D => X"9420B01ACE02152514F80E1249432540090DB900631840814861324C205800CC",
            INIT_RAM_2E => X"39E021B27492909931A1C8844A25108C0C13721B901300213C248A50C02A0C12",
            INIT_RAM_2F => X"4252410A0C64060338A538098F29894C4E1C304B199429270708163090E29484",
            INIT_RAM_30 => X"01FA1A41044024580B018662529139593720025923531BC4CC66C4A18D932610",
            INIT_RAM_31 => X"4210112CA22893408848C1085901E380881A2911132001519CD3B00812828001",
            INIT_RAM_32 => X"DDD1001200D028CDC0C3098A465D1894C0C844D2368C8C1030365A679DA32568",
            INIT_RAM_33 => X"B1A0CA851DCF30CB4641196C209110673998C4EB2599191064C42319B7A42492",
            INIT_RAM_34 => X"99540042C842168966F33448002D76548813128A087890CDA6325010438909B8",
            INIT_RAM_35 => X"A1CCC8441261CD8D2E870257719B0CC0499D00A1386A30084984E06116946645",
            INIT_RAM_36 => X"00434810294E496E4010808884972824CE0488E76CA410B9392313C4220A14D9",
            INIT_RAM_37 => X"D1084089CA098D08CE4366906CDC9106048AE25481048B1CCB3245A231000000",
            INIT_RAM_38 => X"122DCFA46B4502906000101204020000000000B849300088A000AE0D98041094",
            INIT_RAM_39 => X"171ADFFC4926054A20CB493949806AA22A2084482530AC80CE82D8A0CD091867",
            INIT_RAM_3A => X"2203614D83B67244B8C937D5A4480264C05084D41934300A4C9AE4D74AB42B52",
            INIT_RAM_3B => X"17F7763203610810513654E68000050713124810259A0C12D0E4921322890432",
            INIT_RAM_3C => X"76D30678200200BAFE9DDB4D3645889249488F09068F00400830892021864109",
            INIT_RAM_3D => X"55212C410012846909242492A800914256D640516248AAEBFBA966B5835864D0",
            INIT_RAM_3E => X"FA49839821E622580810C8280E480259271829B98319242800100020AA01092A",
            INIT_RAM_3F => X"AAC01801A6C00092D20082506816DB4D12243037924C6800A01600E64A1D27D6"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000200002CFB7BEFFBBFAFFEECAEEFAABFEFBEAFBAFEB00E",
            INIT_RAM_01 => X"040808200440044022010042044108020000000000001C0F0010100000000008",
            INIT_RAM_02 => X"0110010088001002002400140008005001200002002402020002020040800840",
            INIT_RAM_03 => X"F600C104D89DDEE5D59442008460FE002012060BABEBEBFAFEFEBE0000280028",
            INIT_RAM_04 => X"264FB3E5A357BF7D64DDCA53FDCBEEB9ADFABBFEAEDB46DEF0B60BFBF88A8ADE",
            INIT_RAM_05 => X"D4F51120C07ED391D99062292D63AF0473333095951E7965D57CF60CD7A4BC06",
            INIT_RAM_06 => X"24AEF4D4155EA21839D92EFA4DF7A487C6D57D7F9B3CB95A55204208B0FEE51A",
            INIT_RAM_07 => X"AB30FBB396B5A0D3699FC93FD64FFCADBBB7ED9D97BA8BC6BD752CF560CA158A",
            INIT_RAM_08 => X"65B6DCCD453B3CA5F67CBBEFDD96DBECF0D5AFAF1A4C6F5F4FF8F81DFBEE2364",
            INIT_RAM_09 => X"DBFED4C7272637D25E93F0B9A0A838ECA49E0FDDE9022ECBE9FD1DE99E0A23F9",
            INIT_RAM_0A => X"9E1B6FD51A8B84FED5ADCA677F68FB758842D07F4BF77B616582DDC0F3FBC1F5",
            INIT_RAM_0B => X"A3AC8775EBD7FFF946B69FB1A8569FACBEBEEE56539ABEF7AEF0BEBF6F98C44A",
            INIT_RAM_0C => X"1CF1570AC1BE35BC959F74A1F1975F2FA1F19B08D1975E8E38E33A50F0A03577",
            INIT_RAM_0D => X"7D79EBC33CE640443B1BD168F3D5D7BA6AD18C629EB7AC7DC919685500421004",
            INIT_RAM_0E => X"FFDF8B14BDF92D43E4CCD05FCB172C4FAB6DB44ADF6DB6E97BBCCF55180D1C0C",
            INIT_RAM_0F => X"F0C3E3E118FF0E8DF7DF2E6FDC073559AC0D63BA3DF185012CEAD5FF9EFDB944",
            INIT_RAM_10 => X"0F1978C323801120CBB39460C6B06E77F6B57EC387BC5FAFF57076BDDB609C4F",
            INIT_RAM_11 => X"3188F27922432BE1BDAFFC101A980D2000110B45E0107C7E040C05E93E8194C2",
            INIT_RAM_12 => X"0B6A4526C5ED107DAA85143AA01D4540C0202CDBA16CB9A6A92205F28F3278CC",
            INIT_RAM_13 => X"E4F8143F3B64BFED1FFE6DF7E343FFFEB87B877A28CA6B10AB02160BDD55B400",
            INIT_RAM_14 => X"7F09C152667936FF03D3B468477541EAE1EBF5B11112DB164D2652DD610A8A4D",
            INIT_RAM_15 => X"96443E04270B77ADFDC1F2D3911C39BB508D443EC75E3D4A58F06BC8FD7D5104",
            INIT_RAM_16 => X"9CFA7A2006B96191F7356BEF2D963AF7375FF7AFF936DB6B782C4F0F1C525C6F",
            INIT_RAM_17 => X"9BCFEEBE7DC6D2ED75F8ABBF5CDD6E3F59093E7FF56A0FBD9DC979596FD78507",
            INIT_RAM_18 => X"74D35DDD98D64C993266EF9F3B498B5C7DF9E2D7755DDBD14EB4F17C4D7930FA",
            INIT_RAM_19 => X"B2F83EC0D6BC68440A55541EFA62233E79999D75D75D75FFF7267DFF3AFBEFBE",
            INIT_RAM_1A => X"45FF3A776DBDE24933FB4756B5ADA87FF7DF7DE2212F7BDEF54F85FFFF76FDDF",
            INIT_RAM_1B => X"BD6BB5AD6D5556EB45AD6B6A5DDDE660062FBEFBF3FF36E9596596FFEEDECF3F",
            INIT_RAM_1C => X"882F550EE5D7BDEA7EA5ADCFBE8FFB162C476DB6D69553B66F5FBEBD7E96DD2D",
            INIT_RAM_1D => X"5587A967B2DB5F7DDEB63E88CF83BAFEA7FE8B5E3B3C468B1A63C66661C70C98",
            INIT_RAM_1E => X"203DF04769B9B8FA6B19305D81B051D7AF5EAD64D27881BD14B68F8E37C6F9FF",
            INIT_RAM_1F => X"9C7FE033C717B56F6B71FD79D1569D5C7FDBFFFFFFFE3C3C07C1E2E1C04150A4",
            INIT_RAM_20 => X"4516CDCD7D7FDFBD75ADB5B5EF9D5A5F417FEC3BB596F6D7E6EFB32BD3D36874",
            INIT_RAM_21 => X"CD7F1BEDEBDC56DB77BAFD0797F9E98F55BEF1B6FF620019244BF6FB6FF7DC9D",
            INIT_RAM_22 => X"134A061088B59EBD78D9FCFFE4BD1DFB36DFEFFDFEDBD6B7854B7A8B7B27F8E5",
            INIT_RAM_23 => X"5242465D0F0D034082FF37CE7FDD915C681E18DEED0A5BD5B8DF0DFBE0F8E1AB",
            INIT_RAM_24 => X"CF773D05C406D797A947470804FF07803FE0104160ADDD4BF7FFBF7F9C6AAEAC",
            INIT_RAM_25 => X"274942512AF03609A6BC5F11DFCB8B97F86550674E631610421011840FAF06F5",
            INIT_RAM_26 => X"1E68A640C138B9398BE7C5F48A29C12B07C6AAAA215110131543011AA8044244",
            INIT_RAM_27 => X"0096260424B977833878187803838011489C260B8FA888B2E245020A2023C183",
            INIT_RAM_28 => X"30DB6C0002318D57326CCC8BB80389E3494D435C3A010BC1D3420B989C260BBF",
            INIT_RAM_29 => X"C0A7C3DFCB3FC195C01D1BFADD1F2DB703E2A9BB6D5063980EBFADD7E651F98E",
            INIT_RAM_2A => X"9CA7829D307088008994091DCFC810BE68A248AB448F8A91189F859C171F0EFF",
            INIT_RAM_2B => X"6687402424242402334D721212121201D5AF7A0C029C018CA4A704421841308C",
            INIT_RAM_2C => X"5A5A80000000080001B4929900000080FEC0F08430C8010A850EBFFFB7B3B004",
            INIT_RAM_2D => X"E80DC686B7EDFE467815B7C49084809FB4EB2066DFF73BFDF6C06E298BC5E85A",
            INIT_RAM_2E => X"7383877489211F736F15031184C06333A3EB40F2064EB7E5CF893421BCCCB8BD",
            INIT_RAM_2F => X"80648C582191FD68729A63D1265E760B7D60ED36B028C6BC6E6330A7A1CA296B",
            INIT_RAM_30 => X"CDEC411CE18801829AFCEFB58D4126BEE4D6F7F1DEF2FFD266A2ECE499732719",
            INIT_RAM_31 => X"A518083D649208FD9892B083E4431E9C99BE103088D337566ABB884000200020",
            INIT_RAM_32 => X"0AA7607FEC03D1883E492882659B25CE7711DC521D8D92B29DC4F3228F637595",
            INIT_RAM_33 => X"75E63EEE3FF7BEC773B605C148C898C288AD56370B8B0E275EA8E738E090C9A6",
            INIT_RAM_34 => X"8E3E991546B7BDBFC3B2188C0DDAC3CA09950CBEAC2BB783B7E465218431A329",
            INIT_RAM_35 => X"EEC86C4759574BAFD7E8FD9B24B7E2934932DF22B12CE83BF47CAF1CED59523B",
            INIT_RAM_36 => X"6E51355FF08891B81A8777E66CECDEAEF791DBF2C57F7DDFD769EEDBDEBFBDB0",
            INIT_RAM_37 => X"E6F5FDD3962956671CA9DE385BBF6BD25057856B56AF4F91EF2AFF678B4DB6DB",
            INIT_RAM_38 => X"43F91D7D3FCF89F5F8C63580D06835A5B5D45C58D5344444494B2AB89A62211C",
            INIT_RAM_39 => X"861C9CE4C596217A65F66E32839244E4006410347229CDC9C7CB92EE8270740E",
            INIT_RAM_3A => X"A003778F26BA6C10F8EBE5DC3F8506EFE0B1BE59B194E82EED9BFE5B7EEF6F7E",
            INIT_RAM_3B => X"7FDD54CC9E5F19F2D33DD743E0667D3136F2DF5C3FDE5C41BDC1BBB7C19D576F",
            INIT_RAM_3C => X"ADBC139F9FFF2628AD9AB6F1A83E010083823155BEFEEBEE6EA2040CFF158533",
            INIT_RAM_3D => X"D5821C8D666308001000401FFC21E68C02024DD3C005FFFAEAAFC01141F8C056",
            INIT_RAM_3E => X"AFA09468D1E47339F0F7BF716DB6F7F6A6FADF4FC972301C02480491049C21EA",
            INIT_RAM_3F => X"B82491B7348DB649D249B49A6D3492688048624C692A6002001C00001D158764"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FFFFFFFFFFFFFFFFFFFDFFFFCB2DB25B01052BD644517A1110FC410100044FFE",
            INIT_RAM_01 => X"FBF7F7DFFBBFFBBFDDFEFFBDDBBEF7FDFFFFFFFFFFFFE3F0FFEFEFFFFFFFFFF7",
            INIT_RAM_02 => X"FEEFFEFF77FFEFFDFFDBFFEBFFF7FFAFFEDFFFFDFFDBFDFDFFFDFDFFBF7FF7BF",
            INIT_RAM_03 => X"17FD6A32664A570E00E44C98419478F81F0CF86001540155005540FFFFD7FFD7",
            INIT_RAM_04 => X"30405D781130C6602D1011012682CA918024C04AD5048300009146DB0B445188",
            INIT_RAM_05 => X"42DD77038752970B90F0211454D17B8022C970B0C0500B9100010A4800240291",
            INIT_RAM_06 => X"31550A156AA1C0121A92A82D4D962055400000064020820EA2261266D406B404",
            INIT_RAM_07 => X"1008A52396295A8E01B426C004A80300AA01125B8118900340D0BA68F8D6AA33",
            INIT_RAM_08 => X"60B4992050AF34C002582202214936414D4100A0A0D606000CA46D01050BCE97",
            INIT_RAM_09 => X"01685428DAF5A00284488A0D20802080480C07A93BAAC322432150F7BC000039",
            INIT_RAM_0A => X"185E4CE804210300281AB9DD40A04208D6B42A2554A1D0C8C31186B01EA0B725",
            INIT_RAM_0B => X"48C6218488900202C30A0814100208094680011084309A00215B438030538434",
            INIT_RAM_0C => X"E92460853D25697A282955554D54845211A00288540549249088AAAAAA140298",
            INIT_RAM_0D => X"A223232B33155E9112808A3D8940002D42308000910954008D0445044FBDE3FB",
            INIT_RAM_0E => X"000445A9E70456234BBBAA601C81880EBB6DB4E0EE3B6D8452113088A3C7B0F8",
            INIT_RAM_0F => X"2186008A9494E45B2104291A31DF156603B8095016889077042550F60CC7846E",
            INIT_RAM_10 => X"F2AD0035120A0C5496120040102847408C842F813EA81CA1550C1915500A3118",
            INIT_RAM_11 => X"21441B46D1207403100B401A968D4956DB4AD01A15150507B97F7A82F59F98FC",
            INIT_RAM_12 => X"3B3A0B97231FFC6C01CCAF4A5359502E59594400FC0604175ABCF855A02251AA",
            INIT_RAM_13 => X"5B234010D6DB508004110333194084009F08850004108CB5906522DB0C954B35",
            INIT_RAM_14 => X"05D9C150444450522B52B45D56D5406A5549681BBBBA5A5568DAB5B2A6CD5168",
            INIT_RAM_15 => X"82AA828D31448A421A77105064B364400556A2B0AA011A500A0A0038003000A2",
            INIT_RAM_16 => X"7C510822AC282AAA88C0828505C0A0AAE0A1405244345A06C6DAB0A09AE92EA0",
            INIT_RAM_17 => X"311486A829081205154D0EE01320440088B5AF544798BA09551F26082A29521A",
            INIT_RAM_18 => X"F46B555570224489122F4F5065C343D43B553401D77061EC24A25022481490A0",
            INIT_RAM_19 => X"51E622804200287C0BD55408F24001013BBBBDD75D75D77FFF27B55526EBAEBA",
            INIT_RAM_1A => X"01F51241BCED36403368457084200F6AA61861804A54A5294000282545890024",
            INIT_RAM_1B => X"AC42A108400A496844210801C44410A039AEBAEB9555004873CF3C4E2C0C1104",
            INIT_RAM_1C => X"4B0554CA0D406C2B2607150971C9CEB972E0F668077550E2210931D576F40DE8",
            INIT_RAM_1D => X"142C690405214088D6819618650CEB844A5594CBD3E86D76F052D555513AC959",
            INIT_RAM_1E => X"00198080C0C574A551A947535EB888C68D1A28251290A90C45017AF428050500",
            INIT_RAM_1F => X"A0E00027DE1696A06E63409482891226D800000000041C3F0FC1E3C2C0410024",
            INIT_RAM_20 => X"0EC14545555281003C608C0190259F255150AD6A544B09546310556A8AD090C2",
            INIT_RAM_21 => X"B13489B4810F6A4D1804102C44924B2412C0601301A200100236436DB4DB6226",
            INIT_RAM_22 => X"1302054AB2588058B02F40AA061232A5080A82AA00492892062920212074BA8C",
            INIT_RAM_23 => X"120222D0000000857B968EDF52664128300372CFBDFE4B58A4AA1E80038194CC",
            INIT_RAM_24 => X"7A3EAEB1C003681002C5B0F7F800F87FC001EFBE68C0893149081402A8002020",
            INIT_RAM_25 => X"7E4517C8137152BFA42FD000F3EF6A8A6B22AA2E2B71400A0000010A04D6A218",
            INIT_RAM_26 => X"8DFE52B17AF0DD0E773576906C35265A796228A10F396028A9A83A791502E5AB",
            INIT_RAM_27 => X"DD695AAD19EFAEE1FBC8B6366A572CB5A847E59649E25AD60C6357951575ABCD",
            INIT_RAM_28 => X"2FA490000235E75BD387F4E17551EACBBF8B96CB22585710AD96CD7847ACB259",
            INIT_RAM_29 => X"60569004C88300F8782A09AD190E9249F8C28AD249B8A2DC151AD1877FEC3561",
            INIT_RAM_2A => X"AF8240EA3E2E7C00A34F649543E4A06B200C8421180A590E876DA2ACA487234C",
            INIT_RAM_2B => X"0918BFDBDBD9D80284828DEDEDECEC01DDED602F180CA8CAA0C7028404A50AAA",
            INIT_RAM_2C => X"936C77800000000001B4929900000080FEA05A016CA2A4581231400000000005",
            INIT_RAM_2D => X"1424C7541D269C6531301D124843614F91823B025294094B926125595C82056C",
            INIT_RAM_2E => X"29E561322490961925E5D984CA61329489367633B03652510A249210A05D8E24",
            INIT_RAM_2F => X"C252493604C4241338C938149F0DE34DD43424021D8402052109F21090E38489",
            INIT_RAM_30 => X"CFEF00C31E77FC7D5E5BC6FCBC1552123A4350D8E2565BF55591D4404B2ABE8C",
            INIT_RAM_31 => X"DEC5CCE02F96A49403B09CB8D301C36EA085A96D524CCAD929D2033EFF9FBF80",
            INIT_RAM_32 => X"90ABB834A7D188EF4742CAB49499611811147D16A4ACB0DF0447CD28A92B2898",
            INIT_RAM_33 => X"812E1220191756656954C1580284505B1BA1108789D952061C20442176404924",
            INIT_RAM_34 => X"5C152244B098862854B6A006ADFE5A78AA40CD9E2E311BE941D25010409909F7",
            INIT_RAM_35 => X"0ADA8620164BBC0904804016F9F2004ACFF84A283D1477CC4035B6C544944189",
            INIT_RAM_36 => X"0563981031CEC80EC00C442AA7944C2063040843536944037A33B06C621084D5",
            INIT_RAM_37 => X"FF1A9439C2CBAFAA4E056795ECDDB1AFB2669EB19B46AA54D3A2CB8E21A00000",
            INIT_RAM_38 => X"940E07A10302D2C54000052E0D0280010000175A456000000801A89AB0400015",
            INIT_RAM_39 => X"4F5F8D686BAFD0622EDF4F700040720255008790382882E028E2E80DE8203E03",
            INIT_RAM_3A => X"6011628514B026115BDD7557F4F39B5694108E581688779B46CBAE5ACCF6ED67",
            INIT_RAM_3B => X"35757800FE4108DF51E4D6C28048B9F4131F6C1AB11BEF8696409E1B71BB87A6",
            INIT_RAM_3C => X"F4D2175AAD1102208CB9D349F3D0009249499BF1EACEE92322B8A029E5C4C04B",
            INIT_RAM_3D => X"81E50F41005084C909242495540088FF7B7BA0007000EEBFBAFEC1022907F4C0",
            INIT_RAM_3E => X"E6CBA7BC684CCA97583E9300FC9350DF2254C93D0B292A9C00080011003C0A40",
            INIT_RAM_3F => X"FFEDB493FFA49249F6DBFFB6DBEDB7DFB024382721281509E70079C79ED22B36"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"22411114482102912242088926DB4924ABFAAEBFB8BABEEEEBAAABEAFBFEA00B",
            INIT_RAM_01 => X"400080020000800200100800144108922449249249249E9F8911512422491108",
            INIT_RAM_02 => X"8000100800100080020002001000800040020200020040000410001000008000",
            INIT_RAM_03 => X"43AAF55552A97AD52C714A94A55CFE000000000EABFFFEAAAAFFFF8820002000",
            INIT_RAM_04 => X"8ACC9D7A9436AACA86AAAAC64D17E160DCDCD9B260599735B4255555CAA9552D",
            INIT_RAM_05 => X"DEBDF72E9552DE8FF1ED555750557B8551A3B2B16AC567B552AE92AEAAB6B9AA",
            INIT_RAM_06 => X"6560B9555DE8AABA2707A24F532C8AAE962AAAAE5C8A16DCDDAB5AAEAAA9D71F",
            INIT_RAM_07 => X"AB2BBB00A95AE25555AB193260E37C5F41DB648453265D9F97D7BDA8F86D5DAB",
            INIT_RAM_08 => X"8C4924897E7CAAAC56A2AAA4D83249CE916455562AE8F8AAAD54E2D55B6366E0",
            INIT_RAM_09 => X"C8BA2AAE758B5740E313B5D02A208A00EAAEA9B062FBB6C8E2EDC6F7BAAAAA4A",
            INIT_RAM_0A => X"384B5C5108AB979368CAAB751322CBB62D6AE558AB162AAAAAD558C5395DB6ED",
            INIT_RAM_0B => X"8BA6A764CB9BA672973A39C5895639C171566C562AB8AA24ACDB8FBDB983D697",
            INIT_RAM_0C => X"04F5560ACF8CDAD6BC990AAAB1519DB6D454AAAAB000BA28B980855555CAAD64",
            INIT_RAM_0D => X"519E86888AE0A815705D945563901A0D19C94A52963A2A79207172E540000000",
            INIT_RAM_0E => X"A4ED9F3E9CE57DA8ABEFB91BDE3321414492491CAB04926295ECCC77DFAAAA2C",
            INIT_RAM_0F => X"6451CAF07BED9B24DB6CE2659954AAE9F2AB36EA09156E7562AAAE3BBAAC310A",
            INIT_RAM_10 => X"AAAAAAE508D47D55D798B10AC6050B1BA68D7D50BF75555CAAE5662A0BB00C07",
            INIT_RAM_11 => X"5288E4B12A4399EE8EC0B865A812D42DB6D5AAB5CB42AAAEAC5F556A8CAFC55A",
            INIT_RAM_12 => X"54D556AB554EBB5558D353558EC4015EB8B8AACDB576B138E1AAB5555544B3A2",
            INIT_RAM_13 => X"C4ECB9B73124B7B67DB44F7726AAB54CADE64876AAAD534A62E315D47310E45D",
            INIT_RAM_14 => X"5103D6AAAAB1572CAAB54A5D55EAAA95CAAB99C66664A51096256A4E69BBAA96",
            INIT_RAM_15 => X"A85555555555DAC63ED55502EC468CEAB155557CAAAABE5555555573C94AAAAB",
            INIT_RAM_16 => X"C2A2E2AAA94A82AA5D95957150EB355D976CBB2C9142A5B131AD6E5545161C4A",
            INIT_RAM_17 => X"ECEDB1555832B550AAB9C1DD84D572BB654A50ADBB6A6CD943C94DAA85962D6C",
            INIT_RAM_18 => X"0AE8AAAAAAC54A952A522A861DAAA92AABAAE73A28CE9AC15C85C5EC9571255D",
            INIT_RAM_19 => X"EE5832234A4A92A013800516F0AAAAAC4AAAAB2CB2CB2C800552D40011145145",
            INIT_RAM_1A => X"02D8B8726092E5804295B28B5AD5568008A28A2733A318C62AAECEF89F3E7CF9",
            INIT_RAM_1B => X"52B41AD6AAC55495B2D6B5572AAAC710365555557580245A2AAAAAFB94C74CBF",
            INIT_RAM_1C => X"5AAAAB95D2B9D39099C6E3C32C9555AB56B2B0FAA8CAAA9D585CACE669EAC3D5",
            INIT_RAM_1D => X"5D8AD5A0B346ABB431AC508080AB1462244C830773B854C112081575742AA155",
            INIT_RAM_1E => X"A64D994B48AD76DD5D55D566BE1389B162C587575BA8D53940BA6EDC33C67BCF",
            INIT_RAM_1F => X"9119E10F004E20029954D1739B170E5CAED9FFFFFFFC3C0E2FC3E3F3F84252B4",
            INIT_RAM_20 => X"AF9F3AAAAAACF9F9F2D55AAB92102D58B42C55D5CB16472B167E8B5552E3B3B1",
            INIT_RAM_21 => X"CF3659A48B9DE61D24D26AAB16C9AAA655CAE52F2B844901244BD9E79E79E8B8",
            INIT_RAM_22 => X"AF230339C8B95CB962E9F84FCC8C0CF8BA47E4FCBB499793555922DD33318234",
            INIT_RAM_23 => X"5B5556BD5F5F274A9596AD57F34908D1705DC520C0D41DCF184F74D9EE7072BC",
            INIT_RAM_24 => X"6F6687BC6C04914C6AAB8000000000000008000029AFD7C9B9699B14AB557171",
            INIT_RAM_25 => X"7F2E5F4D7BB7F07F9297FDDD9ACF3A0EEB83FF6E7F74773F5AD6D7B76E7CF4AD",
            INIT_RAM_26 => X"D9EE78FDEBF2F16AFF82B7D1CF3873537EB62EBBAFB07628FFD57F7D9FB7F5FF",
            INIT_RAM_27 => X"5D7D5F2E5549B4F5FFE4BB66FF562EB9CDEFFFFE7D235CFB0CAB971FAB9F3E6E",
            INIT_RAM_28 => X"5FDB6FFE64D5EB5DC3AB70EBA7FB3BCBE9AD174DF35D561ABDD70FBDEFFFFE71",
            INIT_RAM_29 => X"B47F71FC5FF76899FE335BADFD5EADB7BBCABBEDB6FEFBDF19BADFD77FE47123",
            INIT_RAM_2A => X"AA085AFF4E8EB634AB9769BFFDEDD695722E8EA32DBE7BBBD77CE3F7FCDD774C",
            INIT_RAM_2B => X"412D3FDBDBD9DBFE00000000000000F15F3BDAA94A3DAB5795F76FCED5AD6AAA",
            INIT_RAM_2C => X"1C7000000000040001B5BA9908080188FFCD3A2D75ABA55ECA5A7FB7FFFBFFFF",
            INIT_RAM_2D => X"4D2E1A1845B6CDAD76916792DAD7E95FD9CCBB777BDE2CE8DB296656A908818F",
            INIT_RAM_2E => X"886F2F32A5B5BE4923D9DAA55AA956A385BE76D3B77E3B65CB25BAB5B6E6DEF4",
            INIT_RAM_2F => X"52D6D75AA41DF44938DD68F09F1DE759D4C5E62E3D8D7F15717B021397E38D7D",
            INIT_RAM_30 => X"8D7B5F58408801001B7BCCECBC5D7E327BC733D9E77B339555D5D4F1D932AE9D",
            INIT_RAM_31 => X"DE16154D6630B9CCDE82F14B555FC77CA32CFD67FB80031DC9C3944080202000",
            INIT_RAM_32 => X"4EFD2376E67B1DEFEE5AEEEAEC192B9C7271C4563C8C95D31C9EDF62AF232739",
            INIT_RAM_33 => X"B5E07AE7BF67A18E53D55C557C1542C72A9CE67F2F991DBE7CEEB39CB27E8492",
            INIT_RAM_34 => X"1DDCFF7C4F9B9EDDC7F63EE3C00E4DDAAF01C5FAF86A30CFB75295B5D48BBB3F",
            INIT_RAM_35 => X"F5D8E377F175FDAF1789BC7A3D5224462BE2B129B8502039C6B466ADF45D7A79",
            INIT_RAM_36 => X"49E2E7EFCDDEDB9EDFD7776EEE8D88A6C654DCCF4C6D5CCB7863B6CDEF3B9ED1",
            INIT_RAM_37 => X"F339CCCBC72B9FEFDE2DE5BBEDCDB39FF736DEF38F6E7E75DF3AC18213892492",
            INIT_RAM_38 => X"55FE9D22572AAAC945AD69561D0A85340555440AE565D5774843BEBAB2EAA53E",
            INIT_RAM_39 => X"1F5FAF7EEBAEFFCF7CBF6B7090D0C55D005555A562AAD78A6B8BE2D6E8721E4E",
            INIT_RAM_3A => X"F013E48FE5F076555BDDBFFFE4F7EE7C9EBBD6F13CA8202E76DFB6F24EB6FFFB",
            INIT_RAM_3B => X"37D5780082EBBD9A7BA67EE7C03FF787B33A6DFBF7B34DD79C65933A73BB9533",
            INIT_RAM_3C => X"249AC66DBBFC4479FE88926B22A489B6DADAABB15EBF54955572ADAE33FC5D7B",
            INIT_RAM_3D => X"7F2B7CD56AF5ADDB5B6D6DAD51AD8FFF7E7EF7FAF24DFABEABAA53977DA776D6",
            INIT_RAM_3E => X"EF8BBFFCF9FFEF78AAF1F93D6F9333DF273A4D1DA30B5501B6D36DA6EFC1ABBF",
            INIT_RAM_3F => X"B8249801B6C00000D249B69349B49268D4ADF32F60086A80080200205EC92F7F"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_basic_kernal
