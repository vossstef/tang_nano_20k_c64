--
--Written by GowinSynthesis
--Tool Version "V1.9.9.01"
--Sat May 11 22:42:12 2024

--Source file index table:
--file0 "\/home/vossstef/Dokumente/tang_nano_20k_c64/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\/home/vossstef/Dokumente/tang_nano_20k_c64/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\/home/vossstef/Gowin_V1.9.9.01_linux/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\/home/vossstef/Gowin_V1.9.9.01_linux/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
vMsGR6KTdoll+1bN+d3MM0FU7G5ZVto0PwGg/ix8M22AIQdoY5eQYmx48dPQNXG2lPykCS7qtH0M
/YxZVwZ1QuqNx819JeIgeYYB5BE7Vjw/4AjWRbR+rGguqk6tq143tKNmYd7KK2C/0UywNWUmmDur
YWaA8mBk40HB3Is/Oi1lCUDGm5tqyDCVOzNcHROeMYSE8U43lhOhvGvreFSSbG3P2WzWqgeAexFy
Jz3X8AZyVkpMjUSkGcNZ+9B8ju5HPgO2QhMYB2rRw0hS4WnveuhxNXNIk0eCIfwlZWz5CL62awHm
6LU6Rn3Dght/VEgWN2CHFHoPe8h+pGbW05ZE0w==

`protect encoding=(enctype="base64", line_length=76, bytes=15360)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
YDfA2VNw9MCcKONamR61c1z+TV8W69ZsNygoxC0xA6uZWyzGHZB2HYZd8gZYWw9BCd8kzMAdoe0X
WG/XvtQsMS1bxeKA61mILSrU7dDd6RcEv/Z9DijuXjI6bBERvVvTU+yhKRpqZQ+ragu7GG7jHh4e
Ki1E/Ib8el3QB6OlDjAhQOuksGrVsqQQenzi8T4NIAkoe5fs4IguKYzY2c0TnuqkReYbkJttuO1P
bxgmRRLRf7Qj9ZcyrorSnlVcGfEAyFzKp2i8MtIXM6Zkges8nXGFGg8uOoDF/PkoT5OU+YxSVqqL
tN9JsRe///Mt76qWP4+MYmPMbDe85FtmxXF7Cj4cZcbIsM2L8QiMYA2Zc7dxVsrzMF+rXf85Erv1
9Bft7op/+E+nBcKxiLvoDW3ZFHvYUwRA44jPsqVQyJYjca9R6ebkzr7DkVrKMxrGDZ9fIWYe26yd
ZBhCfHNmtMrnIcgIpnJYEidv85JwsBeTS/WiGlADLNj85nSNIP7HPu6DdyYY6AsKVznKMmlAlEfJ
s1f4w7HHuaJeCYjL8mCKl2UlF9skpamacsFqq7azBD7fnJPK2f4OyMwxIEWFcsNkSPB39ls7RNpc
FTmh2yMpznmPhJiZ4+RQ+Y+5zW+DV5KjIZHDdCQ/rjtqOapehsQnwwUrPQ1SPLgYm1wPLLS9mspL
Cn1VhDLQoSMDAvy78ilFrp4z8GfUxAeBSLx+cs21Xjc/FNm6JLToKk4aQ6vhcqkU7Lg3Xs/rmGgJ
aCqD8gNk4wyAzysyUXgx/oJVLzFfn/gz3ppOjxQFVI2eO/YKjW50cwNJYArCGmyssq+AwtwmWE9u
50p7F72H5lrUFN3gjJ3/KCiDXhQquhyxnvyxQnEZwR71TosxeSkhyVJKL/ugqVpfWOZo1M6b3RSE
V0PPszwaUDnoUe9SqXyMDj3l4fChJ/T5Zvd+dW1n9SEm+tfMj8/0ApCuhD7yiAAWwKHr8AOln6jA
hnuNDt0SJEuDewohpOwcrzgkeqBexD0THNvqHWTBoCo7S58i/4VBNDLQ92gr00mWPqhUhpSw46JG
KtD40vHcgGA6vx4liOEzWZHO/95jyQiA+u9ISJfQSPAMeMSbuWWn9yAxc+Nbc5/8YGlzP+vMmRjH
E2/tIxW8nlSiiQah06nADUymCQdCd52v8cb4AFeNTXX0ZSmTE0Z8vPK4OOKj8nvdCfvfC2p2r2Oc
vgx4l1f64g3rupJl+AVXAPwRJptZLLY3gimRB8SJs2Hkrz0La8/EYye1Tnil+vZbMYIooIhxhQym
gkOVcBvZEBT1jwcGgYz3/GD83cOhUpLYiXdUTsJQC/vaEXqhTT9NePORRSPUlQ6MfSh8+F/qeBcG
DlmvbyAFFVsJXrxld4ccgD/1R7y19P9CFMARC7fKeTxB1S4joA9T7AGGuRmtc5VIiBbA0z7dzFeg
HEsvGwZRDp7ltcGQtjE3loE/b2wqJQJ8rx+Nhj28PNBm6CcKbVjLkMB6xd2m5RkNtw9kW92s+hxd
iQYS1M+N0Zdp8wIF3E8Rrv2Evz0I+S2RKjJD9Q4M34CxUoZrd2jIkI2+W+BUl1gVZBOfflVvucsh
LMDLX+fY8xmv/vifJegE5qZQaE5XRHPiAOeaQYWDG9EZttPnbzww1TFudgJpjPnCknXPhZ9k2KhU
toYnai+57regxSOLCO8kkNZsCXvRJYKvYQ8DvTmYpzbV67VZT7o8w/3Oqekj3u4/aMZuGPYZW5/c
v6UDy2/Y3ySB3tVHimSheOx3oAoIQyfGGtAhxBNoUgy+28K8dgse72wGhAOeK/k8duiqb1VKM6kI
iMtxqVgfYnrIuFSPZSQKccKWIlHJm8NVwaIIEbMT7uXqFH+uGZhy7kEmFIwbzd/3z+pPYpBRu8DK
Y7nBlRhlX23ptDSVSlT7AGUJpg4OBcljeTSV58yKBCn0/YxcCTCgtokxcx8d6k4IWzCxIbOZp2kr
ibx6EKY8FL9z1eaeM68B9vdKMJofAeME0zI6ha+uWT5zaRs+10T0gTR/nmoQ0wXhNS10GCKj501X
6Zmomm6zJ8x3j/QK19SbN7cYBolP5FOSSZkaGR+sk7Kvm38KiQJHWAEEQPOiNQ8H+qrKou+ST+Ct
6D+gPIncvCi/cTpn+3vr1y5XHb4E2bv9TT84CLCIHVxeNms8S6YGotbW7A8/4zwtl99n1EGYnc/w
KfrzY/S0Dqdl7H5sV7ED862cHl71wo2rAHJ+SwjVSc0+RLCgk2S0yB0sSunH9O97/MsV0Le1uNkT
to3Zuxyrf7p4+bIVW6OnxAp9wjse64PpGDnhJG5qzQ19z86w3cgjN4k+3NKtCVXh9OxQ6JTdjxQj
oAv4xs11qccO23rhUNh+VY8nhXtQeEpr/jdWZqTzlh2VaTs3BRaW/9q7dGM5zhYAc6UY4PHOSC0G
26yECoObIqne9mV2DoGnhDMCz3n+GpluC8ga7YilrmocSU8SgdNr0xyILhxvblqHBn1vB/7x/28n
8muGRqEzO1N4gcSWjaaXetYuBiH+BDCaHFdvjPqj6HtW1NL7uddpmkmy5xBTVoyLH2Obz5sWt5Xl
qwPD4rZsvz8+QPP0yfxS1cgW5Hd2NRCGmS1EqecqOGpcJAFNJQMVPJVBdbmAUbOXoMPrFNXSLvMT
r8tv9ro2hA/fxf9V0N9mK4h7g2mdhISJPH9Bl4X0PXdXawlO3pcCCR60jVR2fi/d4JH5y1DbxOKj
DnUw2KFWyhArNU302HPAc2qNSVsmKdeuEgFs4ij2O1uzaLrknalnc3EtzY5Nt0axPDbHLsrtIC+P
/Vd6Dc5rueelmL7uR1ZWMeX/UM8MDUPplJJqW7QzzQwvG2gD4SyYfpHL8VhzHAR/4tOGOJ1ZWMyd
cF758+O8aQLWjThFtuYHppbLyouIebNUJ3WNeN6C6mmDZRgM1rW1F0x2529LdFVEcYxWeb3EaDU6
SRCWwvcgnrK6rkFJWQ6RORU+yi+TW9vono6gLayrrNRTObGa2UgQCajjvQSEtiEgztDAsC7XLIfd
vOTH2aA/AnqRWt5omSMDNZyNqvmb9WE3lOzrBOCoplwH6to12w0ui2n10YPuBmqKEScc+7qiazYp
dOnicjcVF5qrRv0z2Yka1YNBn6sGsEMjKMno9qR/eqsj6RObnNegHuUZ2q7fRD8H3/RfFTOgB8QX
cj9q+ORYmqUeh4iSjJfSaF3CjXTLosu0QYAmXmq7Y8Hok0/C8tSXrdHGy4TU4urRznnKPYiIozzs
DfavtNqtYy0WIhfMmVTEyBLH9zHriX1UM5o+3gzyzEuwOwYsJIjaz1YKACSYzkWUa78vzyk0h1ws
WMjBu3XLENg3cabiE7UGq4ElqjF7P6wjWWRvX3LVjsyo8kv3S14jwqdgPDHy2NeJRl46sxlIF/xg
pMzdBzxJZJu+IMO4f+D0AAcKxEwNF38wty/gxAUCim/SiBS+NdXKPEZr1rH8oDVJO0ijkc7uHpPX
dB1juTGpk4xJ2heSp1U7yYkPP+zhJJJumasu47ULynXZZIeFzcqkHDm5E6Qu+fpePkQ+f/a+dtmB
PjT55G7IbbKhb0cpSvwEgdJ356fEQF6E7zzmrVFAUr8hko2aKSz7SZ8/4gLT3g/0vl7z+3I8+bA2
jrOoFGx1jYp2N9L0tNjW2P+Yhs6yQgTqPiX2OODP1J1QNObpht7U4pUiNTTJkOxmDto686lWv8JK
Jj5cvPSWhJfivAB4SBEHBnAc/hlkQhWNJa1WBnG/NNWw9vADLBkgme0Ah22NkOtW8B1Sal3ZmTue
jnSyIHqsb4BaWgoq/I/F6Oosh5SD+sa2c/Lfk/kLAabdnnP0FxF7yBqgsD39CM2BqOUe+jLd7Fn+
8TZOVkUquesjSEEC3pCfwMxwBuws3KUM/01p0L/hil636B1vSETgi6AyliGGeNuZLmSxPaqMsc7e
lR4rvSBJ1mTIEEW36FlxQcZ9CVswe56mZlD3Gs77YBhjr/7hx3M+XtIZCtha3zG56/FR0cQL6V1g
ToXz3UngtxltZ82vyn+Bd3nn/kaprTQeRGokPTfsssfbE+MXW0MP6NqQ1uAkgiH46SlJs7E13EFi
yFfP64QdKCqrpuQq01vUFM0waEw/EBE8qwo7j4pohwKW8CGGKXbLZL/1ZGlMo5wqarHSU9ZQNrLk
/1T02JRBqoEwx9hx0JYXfCMd+4yqwURknOvCwc/QedNPMVXipDcU01gLw0RqnFKAndmztymId/tW
4m7leWV0V9f9O2csGgUSYhow1341Hcj5T50pbe3Slc5Ap9QgB7DAPEXgdbklQf8KLcKbGnK20El+
UjIMKroN8gZfGtAj26y/FAfLDWOO6EDZvhonzLiO0F4ZlJ4sOyM9XTkOVE44TFRNDmr+1+26qTM4
/Dj5ReaZILoYSuLs8VAVwpLg7xc+cus/jYlwgJhRl4bbT9xLnGadaoDwXOTNgi97Zpzkj9rkd+n+
fgQDy1MJCcRFwPgvvV/KjmO9YWZFtwLqyZjw4lzjDtg3RYosdlf9N6PhM0S398nrbs1p7M3XzqjO
3S4vglcS/LbnIq6FPT9y7ZCi/F1UFy4oo498qR+ACGYzw9LZ1hyBS+8hjF7e2TmQaVlcTlwrJ5Vk
n7PbW60wnvkrBfOfh3CmQ0XsWinP9a1gYWiX01nrESHfxryJAnVogPOnLl/japg7lCMFsaRxrTk9
8YB+M8ZibVtrl0bl9EZYZlVxVMRYIgCH27jkOUAOKc7902tmlK+bc143yJ+Xv7rYM2shCBY/Yv9n
fu5uEYg56CCgNCtPNnV4FklwM6xpQy3o/eWFRM+yW0IV7zniZGMg/c5fmbIkFk5MF4J8pOhsKMNt
fyh2IAP/UHiiKiaFAr2M4VuzNcg3kUMQOdvzdg7QK5o+TtgVTgtA9YhpzlPY8AnwLthhyo8tVV2v
j89LLdgq7EJVLrqNcx3eHBlQTGY9BE4QpDzKt6mtN0IEqqbhT/lJ3yC98X0zhLlh4qTfayBpSKiO
eYWYCX8H9YEd9UwpqFuRxwFlkuA9M/T4dZLwY8uyC8t2TV9ZTDBmGxT4EQyuIrA3wAsXBe10dYCL
auVN5kmn6LJZaIKUuvYw577fI8v9haHx6+qcE+PqDXoB6585dQPvrJVz9ZdSGd4G2y5AqH6mqwuY
jFtykiMJdgMLM5Va/gVtWHUWOroxrl7VwIg1XpLj6HPNP5vXg/y4Zju85CKz7nBTB6QxWN0w+9gN
6VLIlTOd2WObgTdmai8rIIUirHgTC0C1fmptkkzLM81sRUQbrFESIGb4STUsbPJ/fxQjmO/EC+jW
3UIIbblgE+GpKxUk67RZkFTSjovqcNInW+I05rMrIuV4qp+q55zm0bHwrLAdTnivpoNoDAz3exHC
fYUxshlPI4Ub/JnlGsr6CHR1MfbX6Xap8yeG3YjtZQ7wv2Gi9bF4D+XvjPLVj6lfUMcJqxPD29Kz
acQxuIl2f36IuVC6AwUFzvRYOlI0gPevzxbYyhnQZFwbSWF022NSitwuWpDkNJBwyk7/KwRh1tay
aK8aauw82G29IorUQ6Wf4UmWp8JZ/Z5Y88g51xjTOyFQ+rJ2lqSOtwkfONyxEkzHu5vGlM1uQmT4
kRILyh0gSw7X/AQ5DYbHkP/WR0fpZdIyrE60azouSSzbsIq6vpjyXkRZVI2tkpjqhtAuh+/yIajV
hlij7Ov4rDGC37N+fW5AoYLoKrzUverg2+vI6JSZYRU1tm+rhMRnD5tz+3zrVX89HOoeqRYPKLgq
rPDL1asPX8MWlfmLsS3okM0NFagNVRbZkO5ofesQvq8F1WtmELmMb0dX7AVBw1CBYamSAs6DBsIx
F4Qml2eE1NO9iEpgSrP+LlcykvBepvY6/d/QzXaSkSEDaQ33EemtF9XW/1jkpLZqLuEpl+khfmJc
3qImV+z6cH3tj22D7dPV34O4WbHVhrLI0+l+UHRDbVujkvrqeX4Bbhqh/Mp6sJvSWOPuog5pKBng
IFrV93853EyW00wjPwLq5HUW6j/9dzsTBpGOkPne/qlJ38UrQQB618l7jUuD+VcslrPKa1uKXY2h
5aTw/3fcNv0KA1F6k/DVy84sQNQ3i/cWcU0nu82+T/k10cnhZ6Bu8OduEILfozwqiIrVMOvoBcFT
IV4jkWluNAAEWN0D+bkOeXiUHuQ+lBhjQDrE8OGk49fVpjLPxbBKB2UxorJ+iOu2b+TkvZCnRFRi
fvlxESWs5wnn4DcQVie4jdsas485VFk1tuzVumTHpoCNrFThbF1qPprRwob4Sc15huEW4SNFu0ZK
N5bxTvebWN8plNYnBqP3oU+U9ocSUKII6+f9qlx/GZO2vTIxVmq4XquzQGahoX48dTTK1TdgFoMO
BcASBfTBbawAqMsPbL+Zy9D6JXvnkmWNn+4bJCf0FkNyTAAtncQHjT4Up4qTy/miG5uSafJVb8U6
tJfTlaxCtw/e8jiFT5dMd5dMy72Qoy+DcHolqu27+by16PT6z4injPKizkyPgdoLvLVGemMeEysM
AaQClx8LA1Kepev27/d7aNo+dOnyCYgL5hzmC7ynRt73HH3yRnpZmkP1DwTK6uz4lN/phgQMtBr7
uikTmuCmAGDfAoXgcn0kqEiyhLqt646RBcmNDrdBE1z8QJoH6D8Y/w7fTmLjW5NwmIVXSc3oJfPj
976SQ3tssb4+W9CBkPjWwgQZJtyNnLuMFPIS9JQ20yecpLiaUT2p9Giif5vpLwjVdwvlsie0Rr8E
/Wbn+VRx7Q8dJcNPVgdQvOPF8GiHcNoyIGNG3F4QjQqT5CxU+hvZ37gCxVsHBfd7LtsLTw5zL1G2
eFacFNLB4lu1yd0eGC7YSFy3B8uS6Pyqc/eTAwBb0tcFQXG5dpO4L1sU/kF0QKV2NLV5k5MEa/c/
2M+KhT7w1qPtmWG1pFYidTTO8KEMP7x8mdUSD6pEvB5v+DAhlUKMcw1m5Gg9uDkUsay/NEGtZAWj
hswmD3QM/i1BXh3KgTwUx4hUjNtUONXZ6as5Fb6GIHFPLK6WE607PHcr+Hev3DOmZbZq6RGrCSHW
diytcQQYPDiWBZomi9wUY67q34O0+dNbFl2co6ysATG+sJLNHpNSXE+qx+jU3v8Zsk7dP9B7sO89
V+9rkJSZaW5qGrboD6GoHsO/bosPjkiEzpbHmEJH/Li7TiUIazn+Pe4mzowXCZE0vKE1g0Ot4e0X
yxg3r9MnpFTaxer9Qvww8hVtJo6yaGpy+Dw3Mm8MqyM9rsG18qZsaPDlFBVy8t5NScxYYNsoOBg+
QyWHh4HEn5zH7zcfqBu0zoy085sD8zltYiW/2kMFzW9jdl8ORZX4v7vGdeHDOrrowGmJsUZ1e0PG
mkkAgALcbimY34WXwA+Sv9Ui29cSgMRPxrFRU3LnMYKzmLvsBUthuldVPojyzyYU2Yd1Rqw9Uez7
GzF4aTTM2LJGbcLCbjIvw4KvYe72Z4huK/PyoWtGJVRp5FsoL9VPiEIPK/DHoEvVVXEco563Fv6C
FfTavqCFqBpwLMPnJnXTsbxqdAibBrVCZxNAlZAach2Lo3WyR1fHsFCigSJcynApm8tLgjRtO4jC
grQWW6a6VCsf4hAXUx34+CbrqH1ivW3Drg0Blm6VMo5WGji2nlGFVgi/BjJJ/VLUsmXZ1NuqoiWj
+IfSQhT1US91JaC0SIKzHKL/MX6ISih0Ngn95Fiuvac3T3+iOVPQxffURZddcJhF/6N5Bz3bNUCE
Q7tqiSpnAg0FChhSZRqxsMOBW0/qXZM7Yt8RvL+Py8dRnbQxc1HyuBdTwFzPo7HDqrW9wGm+/uEv
bcZ4lv6Jwq0diCrFyOOffn1xCWl+qSJwiZwJRumvlOXpeoBUR3+gnDaGjfruiSpN4cHBRfdbyuYl
9AhIR9OtyP9oO7GLJHEf3FxHhUJL7Oewa2ZrSwoftyJL1XeN+G6WL22z0V5zbJZEnfjWG0sBiFmG
Vv7I2QhAszZqvyN9o1hQhNADm3WHLbR1Nj1TLeAwvUB4sAYYNpLP7EZoUL2UZPOgwblUhVA9f+68
XQEwgR1Z/YNaME3GjmqHNb8fNZB37YS1+J+QmkT/GcVw0qSkO6xvTelgwKGMyahqH9WieBF5mdnJ
THpb4JCxWoaa+7psNvqYTrHrQja5tEWv0gHBKSJ/BTK5NEb57Cyy0vXa3q7UKmFVmvosTaP5T7gt
XhxqKHlEqldn0kJUi+5Ym4OOCrSEDbJ72GBb15ucUrxG81/t4qk3T1/UB994UOAlGmZ5M22yeam3
zRfsw3GvSEmJJDv9ZH+H+A5hlsYtfzCZyrKQsQ4Q+q2ox96IahbfAps107r4eDVLvCVZmB10fAH9
NMKpck7FKjlD4UuOxH+lGU7mVGcC4guqZYa0YP9aaLGMartUak8EGIm+P9HuubM7ktsI2xoW3LjN
SaIodDEv/SfJAZNufF68m8bFjmnJQMkE9B6eCn8xvkvnx2DqdbyPpj8WNFS6M1txSadVBeaedfmW
m6oimxWjz6G6+7SnBqVmD+741yl1RHVUc1v/g/ltdhhFFgAWGvFbxD2f7Jhvaw7WuseBEhNUtR8C
qfYQb7GLQk1l7Nb50k2RW8iLVmINUrekrzDs+rnRl3A8ycn1uxTagDacG4BNGsjpZfIWwHMYCaJ3
S5URQoYqD2NwKFmMxCkhYPXiBSk5xsvEch8SjUSc8RKVTMQ3iGrnndE0PeujXnC5b0tJnUaprorI
Sz0/jdk1wBP9Cn/UdtIE4/OrOoD7xa3Y0/5vZBZ3G96rFPePB0m85rG2G0Xp82BuH12bxHJasZ6r
fdCJ2Y/LgMoNUUJF33C8bMbHdf2rvT3LPuBZEHpmKCfvu+qrS8uKyCykyCKcllbFZ7ZKgtD7BInN
wI+/dFrc2GkfWn3z4Jifb00prK79fAWERse/gS5H+VCiEORTNcTqf7p4MzxSEB66H8Z36zNq7LZl
LQpkI5n0k3Daym/g76hDHj6zxEhhbG9a1nI5wSXXRt5Vo85DmSvnMysOQ5ZuL/pNM3Cv5454x7MH
3I8z4pUnQKtkbQ1T3ksEQUhSZbxpo9W/p0XC38nesLoy240ZXCUhAnaa0cWLmVSKT+Qzkx/q4Jhu
3Pu/xAgr+SrGG+olHMR9bRcPl8/GuNBMhpDiBbk4lk4NeWYNyrS8CevlrfbrvQN0/bJEv0CnshgL
lL39k9kQ71RfqXyCEbajPeQDH0UqikcQUP/ZKKe3lO8GETfgEHMzK8BQ78HywpdoW8pOoE7/m4Qa
X1/HzjCs9oQvgyuwo4PIk1SKAfvtKGJl1feIb13CU+S0TxX5l9n1eXYOvn9M+OPMsMnS/rPsxNVx
47nNfsiasRwEJl878nK93rr1KA2pqAsm3ECy2CDai2gEl14cPijbMycAa6yuOczy53gFUApm3Psx
zusak1YzG3vUznMhRjvbHzum9/nDVkw4nTFqq8ldQSUEUTuwRfH14VSCMz0kSeUb7WdxUOvK1/52
aab4/CgqaSZkKSL8ukY/8536j6kLNIkPfM2AIPFIM1fT/yLW1ls59dVTuBQOYqR6FHLOknbtiwtL
B7fjbhR3saFpNNyPOjq1gs5GuFZ3J7KZFwvTnkG9hyXFB3UGcxu/ILt9X51fs4/9MYmoIbXvoNNR
xwgzU/6zyXrB0IJS35z5rMoT34siCOVhqhZlvbvTPLyAnbC60NLTHdhlmW0feaaC6tEbUGkhyyTd
V8bkdMm38Zwik/2Vg3gAnoTM5Xw66mk8Ndp1U64oknvs9JC6v5LOFEMXA+u0qp7NrIB4pl1bd5rC
qnDirHrSC8NuOUPPJq51sQ+sFCJU2dKnf1gl07YVedA49yRfTAK1YSaV5fQ2hIwHphQQVQ6QCkzn
dXWUoRcaMCBZijW8knrH0CrRMDPEAPW087AVIZl2vw38O58qZ/QZiOBkEXR7G50n6xgaZOOWgNwm
0sEZtiY5risy+9vKuq7ps5gQyW3huuWZCJ2o0BCJqmsGMDZybkMDUA3L13HI43Bgy3BptRRYcibq
UOnXnalCySiRmyEgBHh2GuWM9+H3lVV9VAh6YsmU8St5/LwWBeWeXe0tCOVCbkROlBAsBMtJujaq
AsM5hnGW5LyCCEe9IGS3v7C6y/B+I3sGQ0bqNj09H38VrJWmyCC7rsAUIxkhg40/YKNI3B5uo4X2
5q6pdF6ZkLbg+pFK8RPjFeuVYO4lwciSplbA2IsbI6L5lJwTFNG6J57wJfR6mEVnOU8stk/4I/Hf
whj92qXbLjKjMpMDxwhNW/Qvcwci8C6e+0T+YTYj5IrFLT5Zgm2jDDm4n+mjuXeZNXuomTt1x4Wn
+ee2SodxR73ltJWEhXK6n11f8kRCNGP5Ss+oe9h3O3ONSj0H97d/mjC23VcGlM8utWuE3CI9HB9B
CvPSS29n4Pn7TM1P6UmmF57wGl8vPb4vyRYppUHW7uHcMnfTTs9WJbqct0YSdwFESM342QG92By+
Qj7mota2Mc0MuwMbNIwUOzWAQnlAdCykk7fI7aV0dDldo9/JLPc5zgaE4c/GPLUXHyEP/bun90FD
9jU7TFQGioCDuRjiSgCnGCR+FgR45aqNU8BStnJY1knO4HiW3c/dksXc6Al7Yd1TnRFO+1ECpxPb
0Qxbqis7beE+e1zKR64GfTzH+cP5ubzXbSmkAgSGSMFBkZN2Yf6AP2WQAQgN5F04yIfPQlWvgRBz
asZZWSkiAHXcKcIer/nOP6JCKxHEPLQJhgJcuad6rx/5dCFTBDBRyIDV+ba84dzsXvTcQajZtYLh
+TzyWTtnCbcF6iBtfsX470zEOsOhqqy1CKOyAr2on7IzerSFBiWJB+/Cwb9dF/61/+DpsoV2ll8c
yCBvvQqGilXXYyEtAaQ/0k4cmxFJFZ8DG3YiveACD8akHuqY6FgRhxpkQ4zp5AZFBmg0mC4QQ9Db
32NPQmtFAX1cuPU0xZh8koTeOCxNY8Ig2WQm396uH/uVVSSVMOGlD8CPByH2pIsgsew7/ACFXV3/
29psWx7HP3x+a6U3NDI7d+ZjQ9l8+/SnWHsDkuNf7CaCsFX9z6aXvKGUbcuyCX8G+BYp8BAhcfS6
O8OqExxy6OUvkrDEnvRlPiJ0Z8Nfnr4kWEuaipdA92unVJ08bKLAVeNXIaeWOGw+3AHemG1WTWXU
1ajqnef61TW9ozL4KqO8iq2RChjXgsV4YqdGS/9FA20YhSAP7mNIPWGQJGB7OJaV7GSDSNwVhvv6
N0yGjLYEwtuNzhH4+XNYIhMpLZ6nIBWkx9LbZcR4Q7rumofGk30cU+54htaizs2clwNlVmA8+o5l
GLyLPhL2pwfLDe2PzIRVq2wR3St10pIDRDKVb8o661Pk5LQqrG/r+aWQCPqtUc/thhXQHRNU+RZD
7X00T+FiubjdOCqrv27IBP7UVKVQ07iQ2B5exsc1jH9kVtbPCLZs/rAH8GvdLQH2y0Mk6XpQLBxq
NK96wZR2GJZo0OTbJgrDA+PMxveeGIqkiQLzlTvPIntlKMhpJdBCpu0VMtAxFHl9c+a0FK0MhD+N
M2Uc9MU8dCLJfpZfLpSCkR/U5VAQa9xhz+XY/yfZbTfNlilcRKrr6Fa4tPYJCqjX7pxSS9rtuvIA
xbd5h6CIjeoI8VgmJzxHm+oF5ebMf2SVq4EHeDUJInFEhS/GkKxsaJB4mWy2GoBVjUqP2M1tJKCG
hIJFethruEsrbSIUonyE1XxhBWyi13UJXMRaWEx38LPr1uVAJQpVZfCdMyfU1zQVrflZkMHwhS6g
YF1gANkHrr9kzViANOX2fc3GrMIQb3ePLmPQEVh153BHm80t4FvNKxTLg1Ju8UABvMztWGAoiJR8
qXdtkDSKAAB7teO0ZAKQCKtogvWvlyrJKseSKX8R76dkpBwKpn/pkjk/z2OHtwWxohkGqf6n6oyc
kNrwhUrF8X1rRhRxYSL7MQ/fWpQ0t1pMQgGmYMKcmaS7yHNj4GmvpkYCGmFeCI1+CZKAOEWaO2lN
QKwIfuwZ86T8VDuFU24eBI5LDQsOZgVfGYypcTijdvuDBLadVQqNI3rYyaFt0Qz3fiWySKGTc7Yk
C6XT9SkdIhgQJNUlrGvC9YdEw+Z59UtH6qoTn7gZo1HeJZ3AMfQ2eqD/Nod07i0ActwEaotxv7yB
TelotYEMUTsC5YAA4QM5PjfwiSkaJNikW0NrpyHo2L8vWDkQ5MvApPj57R9rFT5HvhF/RuJ0Nbtm
OYxw+MXyge2v1hSkdkToSHAtZ2OIXE8RkEj65gTlKwj+CLAtl0yvxZliB3wn7S8DLoEztu584XZ9
+447e/YFoUp69VqXISAZXAlKLlJRNG34Q3E2+GUid3ONrRAcJXa7xruxfrKGDtl2tWEO81YMSzSO
+DCjcBvQuqE4WCmj1zcNUW21kNBjJLVYguywDsPu9CAB1Q0yK4p/vlKxDnwB3sbwSBkevpyI1PT2
nq+8OFuAmfMpdqJbebWfUCBUeKBRcV+gmhO63+7eZOvxdkatQlsHTv2/7vbIrxSz4Z2gvrteCVbZ
xxGr7wzo9CDbsczdxF66M3ihjeHJzRwBmTcXOGKVlug8dfKnUnbnwtdce8hPkos3o67CQjwGI8Z5
U66ftBl6jL6GwCoyc6NWr9Pc4XaeyZoyYFkNRFe/ASxG33lgotwgxvxCYM4aDEGe5TTPeZSmt66d
43s6Ow1wF/I0dYmlT7+A4ADiQX41dXL0r9e7DzoEto3AaT+ZySHW9KHKaTyEy8Nny4IWs/W5u7Rf
UBxJXFhhnSn6Yiar+28NvrCD5hNqPPI21mPEmdqRDPt5SCqU+YJaXYjVcqeld3Nxx6ho0rLBx1hE
1FgLYgor50T2N3YD39qWF3K2/hv7KXRCVyE5an8115gYqOnki5hgkCQ2Okb0QLZRYFsl2MVgkJtC
ZolvfuHw9Qnv9LsgUAAD1ajCt8LZhpPB2/fT2pe+keh8rbT2UgnlkTR5jKmoM2oi2E9Nvg+aBXbR
Nusj5c0iDj6PQDqJ1c2s4l1EsCnakiNQHR+JxkFCiBkae+9gUyEj9wqA3Xc6DZnIBLZlvZmPe4d+
3u3yVTSWTBAJnWYxI/ZvITGhapvQofXsEQIUhIFmIawX4JoqqCPgwHdsqz6qRUJmHLFXD+s5csyP
qiEfTAi89ywtSZ6SUELWTE0HMJbpvB6stJKMfEA/hbmiZAisRF2s4Q7HZgeqIL0PZZCB3IE8XbhL
rJRh7oDfJC5hWHOBeb47pNRylb7bG8XODpTAJnkebXzsTV7SBIzmyL+YA8iUJf7KPMwsbckfcPb7
D5RgWw1jt2r1Ctze7zzexouIcKoEP6EpTh8JfedgKeyCrzdW1ALhojYG6p9cTARJxzjBqKJrguUn
JUZ5RaVRlNzPJQdd86u/NtUEKJxk3niK6+HU81fxiAZi4YB5QWYs9kyn8epc1AV4gVGW+YmHJ/G5
2StxNcWp7+uv2b4z1vG4ATDAo3VC4ieiWdbWkeBv41at7hubvizLSFu3iDAbBYyzjt2Klc/CPWgE
2DZxxkMiNANT1VlY/5jM7aR/drInvk8IP+X1l8wZu6ZozvdxALgtfxgoxHMecMqmpnoN3ETmACFv
ZXrNzCdqdN/+DzHFlGN1hMcB3IBxZ2JNgmMJRnyUKo5I8IzzITDHarhVYupfKpV/HCBw11qVX9/4
Ws+Oj2mwi5S2VaTaTxDMNbhN8SS4UEtOdhv9D/q3FcMf7d3ITrnBxmuCfdDQ2/jPqAEg9Yg0LxK7
p/Obx+46BqdhPq9ZNwAYd86BgTNRHreswFiMUaHVIR2LiRhUrpQ9OT4vEWe0AgCWfypgn4LU3fT2
dVOVlLkzCKXxaL+gRvE3asw1poQpIto00sGenvPqXsQ66kdJYFmi0FXPOA1wVT0iVTShawugWDTV
kAGhjTY3IasrZ/G2WgWQ8g0o8vFuJ/YdpdrF/qSf+QY7tkuKliGpaCWe1U8+h/Plt1YjUzted7Ud
k6dZYDgx4XFnrwJfUHxSsIWBkBxSuwa4H9h3E4WWrruBQRT6pD+6vyeoYTvY9+Lfr1sbSbwXVYU7
V2TQxtwCYL/+NtocrAa2CikrRK6KRkgK7c+JcDlG8oJsUqJiS3o8mEGLA/1yFpDyjrj+VAv/9Unx
VMUj9HyVZYuiaKoEmL3uhmNSXcTXsqqQcYJk7GFhcINqfKruhA2ClGgymZsw4HeNsXOqal9tYTI4
SnxP13AFQVvImfW7smoTRoLgUkIInhFkBN7tp6wY1LJogpk4oJUrfYE8D3bZSvKkZyAsIqCq5jxY
+rrTgacmf+W/S9RvXrvjYn6Hd2A/xl/rlw4+LgFpyGgYfseu0gtX+QcCvHbZriGHuPHkGFHynuR3
FNvPpRzi58w0ahmiTXR743iI4FXJBTYfonPvIIHMllIP/+R8fQlHGNYfTMy4t/UWduV66y91Ud2Q
3W7QqvmYuDzaHUOqaFKc8Z986MHr5ZjO7gJA24AvO80fbZ6o5jORoiOH8aO6EwwDnYvhtagLy7qT
hv2nZUecxKGqeDjOLrKu8e6h/tKeFXtK3wJIlASyvNXI/w6c4zaKU6xY+eC39PaGOOa1vLlYgY/5
ew0c/M5hf7zbSNiG7cBbtMDScECXmBfLf+sd20xe1n762Nbsi6G1TMDR3+i0CKZVLd55OKjKQA04
n9con1W8Bx89Hph3WIRVkVLLM+VahSWcMDFeFBbyoVka8sIB4+eGld9fZnzPFK4teh+9jjss6NGT
Q7Pb7Ol7yx5YGcbuuSmeDC8vau6zDPRzL9UJG5VEqhsYhnf5o35b5RJVwIlj6FEHhIhZaou4/onL
UpXUchIzuA+vwMpppvOnlF3sc+VW24gnXM3+NTtDrWTr/FJzIPyEhWctUkRDk8lunjlQTqyfEyGT
mhI1DVwiBEcpmcQroauXbko+YUgym320+s8Wj97JjgkVuKfLse6ICmCa1pKZfiVhH8ohBJSNhXeb
XbKbX18i6G7dG+XY2ahqzHaXNwoFfSZKeccu40sWppLeSVxprbfkFLJ7zQQTLBDQAfC9i2+EaTS5
TAFzMNbhyVwsub61/mKZN4TnkzBc9f2njSBPMdKwCtKgRO9F/M5AbvIgRKQdUp6Nb2fSC/hlLg9Q
9txF5XvpDKdovMHXO7L/OunYKEzyqhbmA5WXwKtCVv92oI2rIr0FA0r+uZvGxHbJyNq0hP+2I/yZ
kILtd7uxAP8t2ftoqcBKAZcNcgDVwiK69kYpc0p0zphv4lnghNe+23yAgR6lUUCf5yCnF1werXDb
aQeyyV/7YP/uPHmPeg19T01BgjUsH5jYmlKkb1qWnUt4urNYwZMIyHK13+tbNGeVe5TDUJcxESn6
seV1dCR0tBMvVhCLaKTJ3Y7/TfW22qV0/EQhC+0dcVKFT+/F7gYhXaowTYi8wJ7j7Mah/Dbg5Pfz
cv1zbV9ch1pOAcPSjgNhAgvoq/zjIRDM7VsPhD+jv3QY6dIjmxQ2X772rx5gDK5y85T2z5FnxWLc
6CTXhG+tHgnHUpgLdRxybU3uG7dolUCG8FzZGaIzTfw6tloaoSXoO1hAN8CZUoTrgMT3zUHHDQtc
ReXzVd7X8qOSEM/+hDrENXQ/y5L5EGnFnEg8Rk/+RlDjjDsDDoavc0W/X/l0m55WpVlvvB88In5q
Zr2nQylkW/zqccX3fxd0ZLekBwWlmhQGkMiPvxtq2ixkEryPlIfZAT7C+luO0EPQR3MjlbsF04LP
I6iqrEC6TA4JXBecvMem34g927qjf894/z5r7cq5U+/H3zvLnMnxk0I/3I/JfjlY+nCg1RTwFzJa
Axn9tf4bHW4hzLtz+Rf0D2/80FX/wSeEJCrELAsfFbL/zrjJuqT+SmwS1ymmFV8/b77AKJP9JBCb
TA3rMYokUF9i5spm6ZzeAMX7dzFLGVB2XeZ95XsB+k6dk9x3LehrGC2awfz8lRYLfEerF8KDznhD
FzN2H8eT4sLKF8JXsWGmR1E3qoAMdwcBdumTFHX5GxxDzGiyW1n1g3xm1lYs5WsJ0RZ8KdnJ566a
Eo/kf0OS7piecpTV4eDq25fJtxRM678AGs6SlQG13sSzmgeXFSrY0vET4wP5YbxX4SoxzQslQ8tZ
qaVMdZoIvAdk4wJKmlE8fSEe1ddvDdtUecuWRi7LuzQ/2L+lUfzaOG7tqpfm/UN5vyo9nHD+ywdt
heyapHjxzEgf/lOljJo5lFj3O9AoN3eycB4LbVF3gQbV/p6wFIRsVKlLJA6EEX756sE1EsScBjhH
tnxqlVImIviASKMooi5wMFKE+K65vf9hnM0N9pZONz3FVAfd3ObSUF9/MOGNFSTu9l37JKeNfvlH
HEFPdLNUr0DVbUPr9Q3wdtuuDBh2Cw6S0nJm3csEgYF4flkOf3NvDVJ0sxdQSL/KEgXOO0Vkd5sr
TVzJZhCxBsnCIhQSfEIuvz3fT7i2bltzePI7RN8aynjwFTVeftJsbMFvCQf8ctbnYUlCNPFc0hGe
iC5+PvgW8TclC3Q62Uw8hQyBsWwp++35SA5/euHs4ih8k4kq8fXk5ySPeqRrZ9xJjCRH4JiG07fA
hFPtiKqIkgMu1tnHOFW29qL3LYWfmunps2q8Umtu/6sYqnjg/V/NNzn6bPlD1xGL9YBcm/1F5GQD
euPK3aVT4HOQHELGm3i/typX/IISA2TahvMtrzaS/yMW/ozfPDPSe+c1x0aejxKpw/dj9zCtNS/g
xala36h9iqPzD0UJVbHGBA3ZLXfT6NPsCyo2VF8J161bl/v9rftbMMWINzc0Rx5KLbmtSwzNdRUR
SBTpXPJM0VE8t95Ovf3Xx3ZLNahsG74pKWunnZzGiw8ArgFPQfPyJsfZNZHepckJsfxS2Fm+Cae3
FXODHyRdGtVKluKnCvurW8AbScy4tR0b71CZZL6ZmctLrMoS/ahss34xIz1JW1YP24yYzvL8cQOh
WWlxIlrYNky31yWpvDdmVd3SOmJVBab+pjWpUw8JRKDfgG1lbcnEVc/FDGg9ciSWc4YRy8ywU67U
kA3m4lIgygppOQnJmS3ApUvGlmmvK4ehWGzEoqq/0imN0gyrJMOf4T7i4fZLaaEXNLCP5BQtZah8
EO/+NwuOtp+cAT6qBoeeAz0Tb5jQ2b46r4ETBp321rMBuJ31cjPK+f9PRT6cVueqS8JzNDYbpqI3
nD1yNFxwXoGQZNZJ/9S74Jm+jIl2DPENRI34Y9dRlxss3bvbyMvLQu1By6qDAxqjaXnpOaar+yQY
dy2igrdbQ111BtXDnSL5UpdzEdlkLuP6KhTzbkUnQUoENpJ/03e8a7E1oV1hcUQ7Feg1jTCK8J5c
WTK7oj0pShFwgVZfz8j4W7cs78tttwlb0qAQ/B8SAPvizEoZO0TpCi0EgBsICyHYJm1lPAWsVlWx
ZuvIBtzYr5xpv/kCEkneibeCcDd0nTzreY3cbSwiu8tSU3EEOdeQ5G+L7VGjU/He6PadigQeliXk
sZ2cje5gUJidMKEX1eXZ9OFTMzNs5uotvb/X8nA1SwsyGg3iUqcrYfVsg3fimGMc+hsf2nohfNwt
pb6hZmmythkNIi7Lbh/bv5Xim41/s7gwhUwRhde4V0xk7mT4glNJ5XzzFwHTsACaZIR9NfV1EHM6
P4ERsmxY2Bk3slQGeI18z2xPlnKwROP4dgo+AkOzAmvEZDTZaODpMsetlMnqyRrqK1O44RGDAcn9
Y/q5hJk4BHh0XuNakhcVPGsviOcl5/QFut6b9KpMGoiAnW/HlyDASS8BhzWJkfkGBNZcBvDpy6H8
i+638h+RIumhh3jol4XpbP4nQHCBfZFIbXXOotpc//i3kkyqoIcnKiiBFXCdlGkUIazkUVNX5ldg
PXkn5bWyOwBfAquJOc7zkyyl27ettVqSJyG8pMSlT7aUU8x9IQe8/4j1C3KC3ZzfdTrFVC91F25A
Khc8kUwflaY58c5r2EVgvKQMdOHfg9DANXCy+IKBnHCaFNExrMsO+L+TYr+2JMKGt/H/5PYPMce7
MHmQU4CJ9u0Q6fVmvhnRLQe6MRQQSH9f/LK5MOlARpBeUQQ2gsKQ8CZsufffPam7f5QZTM+4Whwv
PLfzTIJ/vL5128WkM3T9t2TCqQnRZyI69v9LV5aswy0XD0/CgSuSvwQLLYIAqtvtoVK0+o0IFU8j
6Edf7r5Vn1wQm5XVRk5ihrY1N5E4uFae6wRh89UJwK2xgaHBvVcFbGhG/pqD/1UlBtupOP5dLzk0
1PUQMJ/NSUwcpdnQB5eK38W5cTwewnPxUoBofa9matZWFixqUwM7pQfcwHneiyFHXUlEpSWFFHIO
WQkj7yi9QRTkTjuSahHPAREVwTH4/JJehErLeNg7dZiOE+zFCt+Orr3M4Z+8mczqEjSrYulOb11F
NK9LpVpG/xtWMLz8/GGmwC/Ra8m/4GG+Zf9etfepFxv4HwJVpxamdjxpdpDqneO34mCABNA8Jhyi
/fZZ+u8hyBT1kEMdswN1V5913tZwy8X/Cuu+uZU4m4bcKmsaTKV2lwzKWbryrXuQOPAN/+H/XfAg
+D8CL7j/nWPp6fePCGjQ/0YoGm8Sfo2XGl56m092YGwBo1TFh1374Aw9jwBUcedVIqYFheo6me3P
bEoxFUoFg51gz/c3yqhuchG53hJVQrWmjNms9LcwHG3c5M20K5HDa/V+GWwADC9GZYTdlJnH1vqa
9i8sgCOITYtDxbyYyanC/WgmMY58T/vEtRXzed7zxnFQ35sAYHVK3xm2tws/hVA/jmiuxWJ+CUhi
sjBg36JoBDHyNzGLezOsxj5eSYbEh8dvG9rIRx83jCpQ06Stzxtg+OrW9U/5yMhVefPRq7Hx2KZu
cpDGi40lBXdTfRMsU3ZdiyuvJnUZizvJ1ShOwqGQOsfgsIyj9NERjPzKavSsRUvoPNGSOkZy6mgo
o6qkSdLQ6wUH5wYzNvO94kUtZXpsDyMkcUeNGnZ4J6OdG5NJWveS20gSedjdvxAZPd+RcYcsJENb
fbHduHXu777ZZtnoo5g1UPaS/YmPvUD42wRFhuhr+i27esBegsRQZJzPYqpj4FKA2ysJqu0pWUWK
6xfLfsdDx1sO5RrQTF7qC+8mLw5auJpuhfAqRc8lGJ9xoRwAHNqdxUZAw0IVNoTBTAfFVI8N54oD
wdeZ6NjMI5ZEFEb4Um2IAHzIZXXERl97XWzrHHxNxolm8T8qC5HiUHc5e+V/2v0iAESMrrzXgagm
BOeCuhOi1SNSVN3bHXOhnqoq1WGR1dpEBEngoPiKXmFJjprHmvOEayM1AZCYiJtsWLDOtR4snzXF
jcCDvycHikDSVHIv5DE/nN13Ltm1wSO9augTUp0ljwRZssvY7McfNlPmxwknpMsGphFw/I+4nBN2
i5/15gxaRXsS5NXvSYJu8RmiA6beWRbn5SGoj0Wfjv5O2++qVaMUnHv6FIE0yeujwxJcV4Ikot6H
suS9XVDBpqVU6JxD1hnuRt36i7G4LjQ+18WxVMrKh/mYj/pGzWbIhC0tspXjY96EoiEuBZyMif3G
Xyjo4qU8GbgdBs+3vYjEPvFpTC7YXd3cdNTDPjRaDkU7Qgbgg9rXNlfe2E10BrP6Tv2jEghNIbNE
CA1Q1oa1/3uYg6McZJUWN08nSFMT651OI6x8SLhrPlhBVTWzXga5d9etk0v/akO7+KmtgQjPguj3
Q3aO+yKQd/XlyrAmb27rVab3W/6krmQBSS7pKkoW6XLGiSQuc7T7MsWspZBdPvJ4Lk55xm1lKY4D
NQ7olJb/cKw4k5oaDNNWoPRpJ5kaGlbS17m6Zr1ZgFvCu8SmSVzoLTQMuWIt5fGSw0Gl+DmWxxZ0
ge7cTBa1T9EeuFOTP1aoqnpA27MSmtH1CdVx+pkkrSY1wWk/r/Rk076vmQmXDZOUdpAdzQ42ArvK
j0slExw5JLGag9nHLifXOwtWsp83+n2a+KlWYTA0OdK6GX9bC7Urv/NTDHkg3iBkGc0/ehjX25qL
9FDVW/EJ5mJ9mmMpAD56m7K+LCaR+7zkMR0wSl5snFtC8S2TZuS0VxlDQO3HlVCScZYY1BfsIhHK
ikAEWi4HTtNVx98Jmef9GtvOH4bO/aWPj6pqZiizC1ZTCC6vfT5Z687VYK1AgpWYfnHldlGIs1rg
bYHvo0aoESuu/Zb4h60PG3vbpm3cC7d3B1HlWbf5Ep6YZHAJyUb1fJ4VnTvLwsS7g1HbBObJNogY
ZvSQt62TtZ2xWxEmK1Q8LG+zjwKJ6FFdAaOOsjImeEMRST9uLp6q9JCFXgUo50Om9kxwKDMNxZl7
Ht5TEwq3otc5BisNowqmvMiHC2sSs/6DnyCd+izNXhYdbtzOjoD10Yc+bteRNdUrk6pXVnUQjFTD
XcBhZq1T377wESbadn7wb01CoAgH/E/ua9DzWWeNJ/1405EJGpNQ47PHSOodJDYiyV1OnIzrqk79
qlJs8SmHQXbAN4u0WKNMoDGI/lp3ose3l/Ki
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity FIFO_SC_HS_Top is
port(
  Data :  in std_logic_vector(7 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(7 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end FIFO_SC_HS_Top;
architecture beh of FIFO_SC_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo_sc_hs.FIFO_SC_HS_Top\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(7 downto 0);
  Full: out std_logic;
  Empty: out std_logic;
  Q : out std_logic_vector(7 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.FIFO_SC_HS_Top\
port map(
  Clk => Clk,
  Reset => Reset,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(7 downto 0) => Data(7 downto 0),
  Full => NN_0,
  Empty => NN,
  Q(7 downto 0) => Q(7 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
